`include "SIMON_defintions.svh"

module test_SIMON_topPKT_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define	PKT_MAX 1259
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;

        inPKT[0]        = 80'hE0001918111009080100;
        inPKT[1]        = 80'hC0016565687765656877;
        inPKT[2]        = 80'hC002446F6E6563207365;
        inPKT[3]        = 80'hC00364206E756C6C6120;
        inPKT[4]        = 80'hC00475726E612E204E75;
        inPKT[5]        = 80'hC0056C6C616D20616320;
        inPKT[6]        = 80'hC0066461706962757320;
        inPKT[7]        = 80'hC0076C6967756C612E20;
        inPKT[8]        = 80'hC008436C617373206170;
        inPKT[9]        = 80'hC00974656E7420746163;
        inPKT[10]       = 80'hC00A69746920736F6369;
        inPKT[11]       = 80'hC00B6F73717520616420;
        inPKT[12]       = 80'hC00C6C69746F72612074;
        inPKT[13]       = 80'hC00D6F727175656E7420;
        inPKT[14]       = 80'hC00E70657220636F6E75;
        inPKT[15]       = 80'hC00F626961206E6F7374;
        inPKT[16]       = 80'hC01072612C2070657220;
        inPKT[17]       = 80'hC011696E636570746F73;
        inPKT[18]       = 80'hC0122068696D656E6165;
        inPKT[19]       = 80'hC0136F732E2053757370;
        inPKT[20]       = 80'hC014656E646973736520;
        inPKT[21]       = 80'hC0156665726D656E7475;
        inPKT[22]       = 80'hC0166D20707572757320;
        inPKT[23]       = 80'hC0176E6F6E206E756E63;
        inPKT[24]       = 80'hC0182066617563696275;
        inPKT[25]       = 80'hC019732C20696E20706C;
        inPKT[26]       = 80'hC01A6163657261742061;
        inPKT[27]       = 80'hC01B6E746520636F6E67;
        inPKT[28]       = 80'hC01C75652E204D617572;
        inPKT[29]       = 80'hC01D697320696163756C;
        inPKT[30]       = 80'hC01E6973207574206D61;
        inPKT[31]       = 80'hC01F676E612076656C20;
        inPKT[32]       = 80'hC020646170696275732E;
        inPKT[33]       = 80'hC0212043757261626974;
        inPKT[34]       = 80'hC0227572207361676974;
        inPKT[35]       = 80'hC02374697320616E7465;
        inPKT[36]       = 80'hC024206D61676E612E20;
        inPKT[37]       = 80'hC025496E2074656D706F;
        inPKT[38]       = 80'hC02672206C6F72656D20;
        inPKT[39]       = 80'hC0276C6F72656D2C206E;
        inPKT[40]       = 80'hC0286F6E206D61747469;
        inPKT[41]       = 80'hC0297320617263752076;
        inPKT[42]       = 80'hC02A6976657272612065;
        inPKT[43]       = 80'hC02B752E20436C617373;
        inPKT[44]       = 80'hC02C20617074656E7420;
        inPKT[45]       = 80'hC02D7461636974692073;
        inPKT[46]       = 80'hC02E6F63696F73717520;
        inPKT[47]       = 80'hC02F6164206C69746F72;
        inPKT[48]       = 80'hC0306120746F72717565;
        inPKT[49]       = 80'hC0316E74207065722063;
        inPKT[50]       = 80'hC0326F6E75626961206E;
        inPKT[51]       = 80'hC0336F737472612C2070;
        inPKT[52]       = 80'hC034657220696E636570;
        inPKT[53]       = 80'hC035746F732068696D65;
        inPKT[54]       = 80'hC0366E61656F732E2056;
        inPKT[55]       = 80'hC0376573746962756C75;
        inPKT[56]       = 80'hC0386D2073656420616C;
        inPKT[57]       = 80'hC039697175616D206C65;
        inPKT[58]       = 80'hC03A637475732C207075;
        inPKT[59]       = 80'hC03B6C76696E61722061;
        inPKT[60]       = 80'hC03C6C697175616D206C;
        inPKT[61]       = 80'hC03D616375732E204D6F;
        inPKT[62]       = 80'hC03E7262692061726375;
        inPKT[63]       = 80'hC03F20697073756D2C20;
        inPKT[64]       = 80'hC0407363656C65726973;
        inPKT[65]       = 80'hC041717565206E6F6E20;
        inPKT[66]       = 80'hC0427075727573207574;
        inPKT[67]       = 80'hC0432C20706C61636572;
        inPKT[68]       = 80'hC0446174206665726D65;
        inPKT[69]       = 80'hC0456E74756D206C656F;
        inPKT[70]       = 80'hC0462E20517569737175;
        inPKT[71]       = 80'hC0476520617563746F72;
        inPKT[72]       = 80'hC0482073697420616D65;
        inPKT[73]       = 80'hC0497420617263752075;
        inPKT[74]       = 80'hC04A74206D616C657375;
        inPKT[75]       = 80'hC04B6164612E20557420;
        inPKT[76]       = 80'hC04C74696E636964756E;
        inPKT[77]       = 80'hC04D74206D61676E6120;
        inPKT[78]       = 80'hC04E72686F6E63757320;
        inPKT[79]       = 80'hC04F6772617669646120;
        inPKT[80]       = 80'hC050626C616E6469742E;
        inPKT[81]       = 80'hC0510D0A0D0A446F6E65;
        inPKT[82]       = 80'hC0526320696E20646961;
        inPKT[83]       = 80'hC0536D206E756E632E20;
        inPKT[84]       = 80'hC05453757370656E6469;
        inPKT[85]       = 80'hC0557373652076656C20;
        inPKT[86]       = 80'hC056646F6C6F72207669;
        inPKT[87]       = 80'hC057746165206D617572;
        inPKT[88]       = 80'hC05869732070656C6C65;
        inPKT[89]       = 80'hC0596E74657371756520;
        inPKT[90]       = 80'hC05A706C616365726174;
        inPKT[91]       = 80'hC05B207574206574206D;
        inPKT[92]       = 80'hC05C692E205072616573;
        inPKT[93]       = 80'hC05D656E742076656C20;
        inPKT[94]       = 80'hC05E656E696D20696420;
        inPKT[95]       = 80'hC05F6A7573746F206D61;
        inPKT[96]       = 80'hC0606C65737561646120;
        inPKT[97]       = 80'hC061756C6C616D636F72;
        inPKT[98]       = 80'hC0627065722E204D6F72;
        inPKT[99]       = 80'hC06362692068656E6472;
        inPKT[100]      = 80'hC0646572697420666572;
        inPKT[101]      = 80'hC0656D656E74756D2065;
        inPKT[102]      = 80'hC0666E696D2073697420;
        inPKT[103]      = 80'hC067616D6574206C6163;
        inPKT[104]      = 80'hC068696E69612E204165;
        inPKT[105]      = 80'hC0696E65616E2073656D;
        inPKT[106]      = 80'hC06A206475692C206661;
        inPKT[107]      = 80'hC06B7563696275732075;
        inPKT[108]      = 80'hC06C74206C6967756C61;
        inPKT[109]      = 80'hC06D2073697420616D65;
        inPKT[110]      = 80'hC06E742C20696D706572;
        inPKT[111]      = 80'hC06F6469657420636F6D;
        inPKT[112]      = 80'hC0706D6F646F206E6973;
        inPKT[113]      = 80'hC0716C2E205175697371;
        inPKT[114]      = 80'hC0727565206F64696F20;
        inPKT[115]      = 80'hC0736D61757269732C20;
        inPKT[116]      = 80'hC074766573746962756C;
        inPKT[117]      = 80'hC075756D20616320696E;
        inPKT[118]      = 80'hC07674657264756D2069;
        inPKT[119]      = 80'hC077642C206567657374;
        inPKT[120]      = 80'hC0786173206E6F6E2064;
        inPKT[121]      = 80'hC07975692E204E756E63;
        inPKT[122]      = 80'hC07A2065666669636974;
        inPKT[123]      = 80'hC07B75722C2072697375;
        inPKT[124]      = 80'hC07C7320656765742076;
        inPKT[125]      = 80'hC07D656E656E61746973;
        inPKT[126]      = 80'hC07E2076656E656E6174;
        inPKT[127]      = 80'hC07F69732C2065726F73;
        inPKT[128]      = 80'hC080206E697369206961;
        inPKT[129]      = 80'hC08163756C6973206E75;
        inPKT[130]      = 80'hC0826C6C612C20696E20;
        inPKT[131]      = 80'hC08376756C7075746174;
        inPKT[132]      = 80'hC084652075726E61206F;
        inPKT[133]      = 80'hC08564696F2065676574;
        inPKT[134]      = 80'hC086206C616375732E20;
        inPKT[135]      = 80'hC087566976616D757320;
        inPKT[136]      = 80'hC088636F6E7365717561;
        inPKT[137]      = 80'hC0897420766172697573;
        inPKT[138]      = 80'hC08A206E756C6C612C20;
        inPKT[139]      = 80'hC08B6163206469676E69;
        inPKT[140]      = 80'hC08C7373696D206C6563;
        inPKT[141]      = 80'hC08D7475732E0D0A0D0A;
        inPKT[142]      = 80'hC08E446F6E6563206961;
        inPKT[143]      = 80'hC08F63756C6973206E75;
        inPKT[144]      = 80'hC0906E6320696E206C6F;
        inPKT[145]      = 80'hC09172656D2073616769;
        inPKT[146]      = 80'hC092747469732C206575;
        inPKT[147]      = 80'hC0932073616769747469;
        inPKT[148]      = 80'hC094732074656C6C7573;
        inPKT[149]      = 80'hC0952073616769747469;
        inPKT[150]      = 80'hC096732E205665737469;
        inPKT[151]      = 80'hC09762756C756D206C69;
        inPKT[152]      = 80'hC0986265726F206D6175;
        inPKT[153]      = 80'hC0997269732C20766F6C;
        inPKT[154]      = 80'hC09A7574706174206120;
        inPKT[155]      = 80'hC09B6E756E63206E6563;
        inPKT[156]      = 80'hC09C2C20616C69717561;
        inPKT[157]      = 80'hC09D6D20706861726574;
        inPKT[158]      = 80'hC09E726120657261742E;
        inPKT[159]      = 80'hC09F20566976616D7573;
        inPKT[160]      = 80'hC0A0206175677565206A;
        inPKT[161]      = 80'hC0A17573746F2C206772;
        inPKT[162]      = 80'hC0A26176696461206575;
        inPKT[163]      = 80'hC0A320756C6C616D636F;
        inPKT[164]      = 80'hC0A472706572206E6563;
        inPKT[165]      = 80'hC0A52C20637572737573;
        inPKT[166]      = 80'hC0A6206174206C6F7265;
        inPKT[167]      = 80'hC0A76D2E204475697320;
        inPKT[168]      = 80'hC0A86C75637475732065;
        inPKT[169]      = 80'hC0A97374206964206E69;
        inPKT[170]      = 80'hC0AA62682074696E6369;
        inPKT[171]      = 80'hC0AB64756E742C207574;
        inPKT[172]      = 80'hC0AC20636F6E73656374;
        inPKT[173]      = 80'hC0AD657475722065726F;
        inPKT[174]      = 80'hC0AE7320666575676961;
        inPKT[175]      = 80'hC0AF742E2041656E6561;
        inPKT[176]      = 80'hC0B06E2073656D706572;
        inPKT[177]      = 80'hC0B120636F6E67756520;
        inPKT[178]      = 80'hC0B26C65637475732C20;
        inPKT[179]      = 80'hC0B36E6563206665726D;
        inPKT[180]      = 80'hC0B4656E74756D206C65;
        inPKT[181]      = 80'hC0B56F20636F6E677565;
        inPKT[182]      = 80'hC0B620717569732E204D;
        inPKT[183]      = 80'hC0B76F7262692076756C;
        inPKT[184]      = 80'hC0B87075746174652069;
        inPKT[185]      = 80'hC0B96D70657264696574;
        inPKT[186]      = 80'hC0BA2075726E61207574;
        inPKT[187]      = 80'hC0BB2074696E63696475;
        inPKT[188]      = 80'hC0BC6E742E204D616563;
        inPKT[189]      = 80'hC0BD656E617320657520;
        inPKT[190]      = 80'hC0BE6D69206E756C6C61;
        inPKT[191]      = 80'hC0BF2E20457469616D20;
        inPKT[192]      = 80'hC0C0656C697420697073;
        inPKT[193]      = 80'hC0C1756D2C20706C6163;
        inPKT[194]      = 80'hC0C26572617420656765;
        inPKT[195]      = 80'hC0C37420706861726574;
        inPKT[196]      = 80'hC0C47261206E65632C20;
        inPKT[197]      = 80'hC0C5617563746F722061;
        inPKT[198]      = 80'hC0C6207175616D2E2049;
        inPKT[199]      = 80'hC0C76E2076656C206961;
        inPKT[200]      = 80'hC0C863756C6973206F64;
        inPKT[201]      = 80'hC0C9696F2E204E756C6C;
        inPKT[202]      = 80'hC0CA616D2076656C2064;
        inPKT[203]      = 80'hC0CB69676E697373696D;
        inPKT[204]      = 80'hC0CC206E756E632C2076;
        inPKT[205]      = 80'hC0CD6974616520636F6E;
        inPKT[206]      = 80'hC0CE7365717561742074;
        inPKT[207]      = 80'hC0CF75727069732E2043;
        inPKT[208]      = 80'hC0D07572616269747572;
        inPKT[209]      = 80'hC0D1206575206D692064;
        inPKT[210]      = 80'hC0D269676E697373696D;
        inPKT[211]      = 80'hC0D32C206D6F6C6C6973;
        inPKT[212]      = 80'hC0D42070757275732061;
        inPKT[213]      = 80'hC0D5632C20657569736D;
        inPKT[214]      = 80'hC0D66F64206C69626572;
        inPKT[215]      = 80'hC0D76F2E2050656C6C65;
        inPKT[216]      = 80'hC0D86E74657371756520;
        inPKT[217]      = 80'hC0D96E756E6320656E69;
        inPKT[218]      = 80'hC0DA6D2C20636F6E6469;
        inPKT[219]      = 80'hC0DB6D656E74756D2076;
        inPKT[220]      = 80'hC0DC656C2065726F7320;
        inPKT[221]      = 80'hC0DD65752C20696D7065;
        inPKT[222]      = 80'hC0DE726469657420696D;
        inPKT[223]      = 80'hC0DF7065726469657420;
        inPKT[224]      = 80'hC0E070757275732E0D0A;
        inPKT[225]      = 80'hC0E10D0A437261732070;
        inPKT[226]      = 80'hC0E2656C6C656E746573;
        inPKT[227]      = 80'hC0E3717565206D617572;
        inPKT[228]      = 80'hC0E46973207175697320;
        inPKT[229]      = 80'hC0E56D61757269732073;
        inPKT[230]      = 80'hC0E663656C6572697371;
        inPKT[231]      = 80'hC0E7756520756C747269;
        inPKT[232]      = 80'hC0E86369657320736974;
        inPKT[233]      = 80'hC0E920616D657420696E;
        inPKT[234]      = 80'hC0EA206C616375732E20;
        inPKT[235]      = 80'hC0EB4D6175726973206C;
        inPKT[236]      = 80'hC0EC6F626F7274697320;
        inPKT[237]      = 80'hC0ED7269737573207175;
        inPKT[238]      = 80'hC0EE697320657820756C;
        inPKT[239]      = 80'hC0EF7472696365732063;
        inPKT[240]      = 80'hC0F06F6E736563746574;
        inPKT[241]      = 80'hC0F175722E204E756C6C;
        inPKT[242]      = 80'hC0F261206D6174746973;
        inPKT[243]      = 80'hC0F3206E696268207369;
        inPKT[244]      = 80'hC0F47420616D65742064;
        inPKT[245]      = 80'hC0F569616D2072686F6E;
        inPKT[246]      = 80'hC0F66375732C20736974;
        inPKT[247]      = 80'hC0F720616D6574207665;
        inPKT[248]      = 80'hC0F873746962756C756D;
        inPKT[249]      = 80'hC0F920746F72746F7220;
        inPKT[250]      = 80'hC0FA7072657469756D2E;
        inPKT[251]      = 80'hC0FB204E756C6C612076;
        inPKT[252]      = 80'hC0FC656E656E61746973;
        inPKT[253]      = 80'hC0FD206469616D206665;
        inPKT[254]      = 80'hC0FE6C69732C20657420;
        inPKT[255]      = 80'hC0FF6665756769617420;
        inPKT[256]      = 80'hC000746F72746F722074;
        inPKT[257]      = 80'hC0017269737469717565;
        inPKT[258]      = 80'hC0022076697461652E20;
        inPKT[259]      = 80'hC0034E756C6C61206672;
        inPKT[260]      = 80'hC004696E67696C6C6120;
        inPKT[261]      = 80'hC005646F6C6F72206D69;
        inPKT[262]      = 80'hC0062C20757420636F6E;
        inPKT[263]      = 80'hC00776616C6C69732065;
        inPKT[264]      = 80'hC0086C697420756C7472;
        inPKT[265]      = 80'hC0096963657320612E20;
        inPKT[266]      = 80'hC00A44756973206C6F62;
        inPKT[267]      = 80'hC00B6F7274697320706F;
        inPKT[268]      = 80'hC00C72747469746F7220;
        inPKT[269]      = 80'hC00D636F6E76616C6C69;
        inPKT[270]      = 80'hC00E732E20457469616D;
        inPKT[271]      = 80'hC00F2065726174206A75;
        inPKT[272]      = 80'hC01073746F2C20706F73;
        inPKT[273]      = 80'hC0117565726520717569;
        inPKT[274]      = 80'hC0127320706F73756572;
        inPKT[275]      = 80'hC013652061632C20636F;
        inPKT[276]      = 80'hC0146D6D6F646F207669;
        inPKT[277]      = 80'hC015746165206D617373;
        inPKT[278]      = 80'hC016612E204375726162;
        inPKT[279]      = 80'hC0176974757220746F72;
        inPKT[280]      = 80'hC018746F722074757270;
        inPKT[281]      = 80'hC01969732C2074696E63;
        inPKT[282]      = 80'hC01A6964756E74206964;
        inPKT[283]      = 80'hC01B206672696E67696C;
        inPKT[284]      = 80'hC01C6C612065752C2076;
        inPKT[285]      = 80'hC01D6F6C757470617420;
        inPKT[286]      = 80'hC01E6174206C6967756C;
        inPKT[287]      = 80'hC01F612E205365642073;
        inPKT[288]      = 80'hC0206167697474697320;
        inPKT[289]      = 80'hC021617420697073756D;
        inPKT[290]      = 80'hC0222061742062696265;
        inPKT[291]      = 80'hC0236E64756D2E20416C;
        inPKT[292]      = 80'hC024697175616D206567;
        inPKT[293]      = 80'hC025657420706F727461;
        inPKT[294]      = 80'hC0262076656C69742E20;
        inPKT[295]      = 80'hC0274E756E6320616363;
        inPKT[296]      = 80'hC028756D73616E207072;
        inPKT[297]      = 80'hC029657469756D206D61;
        inPKT[298]      = 80'hC02A676E612C2070656C;
        inPKT[299]      = 80'hC02B6C656E7465737175;
        inPKT[300]      = 80'hC02C652072686F6E6375;
        inPKT[301]      = 80'hC02D732065782074696E;
        inPKT[302]      = 80'hC02E636964756E742076;
        inPKT[303]      = 80'hC02F697461652E20446F;
        inPKT[304]      = 80'hC0306E6563207574206E;
        inPKT[305]      = 80'hC03169626820616E7465;
        inPKT[306]      = 80'hC0322E20437572616269;
        inPKT[307]      = 80'hC03374757220656C656D;
        inPKT[308]      = 80'hC034656E74756D2C2071;
        inPKT[309]      = 80'hC03575616D2061632073;
        inPKT[310]      = 80'hC036656D706572206C75;
        inPKT[311]      = 80'hC037637475732C20616E;
        inPKT[312]      = 80'hC0387465206578206567;
        inPKT[313]      = 80'hC0396573746173207269;
        inPKT[314]      = 80'hC03A7375732C20616320;
        inPKT[315]      = 80'hC03B6D6178696D757320;
        inPKT[316]      = 80'hC03C7175616D20717561;
        inPKT[317]      = 80'hC03D6D20766974616520;
        inPKT[318]      = 80'hC03E656C69742E204D6F;
        inPKT[319]      = 80'hC03F7262692065676574;
        inPKT[320]      = 80'hC0402061726375207369;
        inPKT[321]      = 80'hC0417420616D6574206C;
        inPKT[322]      = 80'hC0426967756C6120706F;
        inPKT[323]      = 80'hC043727461206D617474;
        inPKT[324]      = 80'hC04469732E204D616563;
        inPKT[325]      = 80'hC045656E61732074696E;
        inPKT[326]      = 80'hC046636964756E742061;
        inPKT[327]      = 80'hC0477567756520646170;
        inPKT[328]      = 80'hC0486962757320657374;
        inPKT[329]      = 80'hC04920756C6C616D636F;
        inPKT[330]      = 80'hC04A7270657220656765;
        inPKT[331]      = 80'hC04B737461732E0D0A0D;
        inPKT[332]      = 80'hC04C0A4D6F7262692065;
        inPKT[333]      = 80'hC04D7569736D6F642066;
        inPKT[334]      = 80'hC04E6575676961742064;
        inPKT[335]      = 80'hC04F6F6C6F722076656C;
        inPKT[336]      = 80'hC0502064617069627573;
        inPKT[337]      = 80'hC0512E204D616563656E;
        inPKT[338]      = 80'hC0526173207361676974;
        inPKT[339]      = 80'hC0537469732065666669;
        inPKT[340]      = 80'hC0546369747572206572;
        inPKT[341]      = 80'hC0556F732C206964206C;
        inPKT[342]      = 80'hC0566F626F7274697320;
        inPKT[343]      = 80'hC057616E746520736365;
        inPKT[344]      = 80'hC0586C65726973717565;
        inPKT[345]      = 80'hC0592072686F6E637573;
        inPKT[346]      = 80'hC05A2E20496E20616C69;
        inPKT[347]      = 80'hC05B7175616D2C206572;
        inPKT[348]      = 80'hC05C6174206D61747469;
        inPKT[349]      = 80'hC05D7320706C61636572;
        inPKT[350]      = 80'hC05E6174206567657374;
        inPKT[351]      = 80'hC05F61732C20746F7274;
        inPKT[352]      = 80'hC0606F7220746F72746F;
        inPKT[353]      = 80'hC0617220626C616E6469;
        inPKT[354]      = 80'hC062742073656D2C206E;
        inPKT[355]      = 80'hC063656320636F6E7661;
        inPKT[356]      = 80'hC0646C6C69732075726E;
        inPKT[357]      = 80'hC0656120656C69742065;
        inPKT[358]      = 80'hC06674206F64696F2E20;
        inPKT[359]      = 80'hC067566573746962756C;
        inPKT[360]      = 80'hC068756D206964206C65;
        inPKT[361]      = 80'hC0696F2066656C69732E;
        inPKT[362]      = 80'hC06A204E756E6320706F;
        inPKT[363]      = 80'hC06B72747469746F7220;
        inPKT[364]      = 80'hC06C617563746F722071;
        inPKT[365]      = 80'hC06D75616D2C20656C65;
        inPKT[366]      = 80'hC06E6D656E74756D2076;
        inPKT[367]      = 80'hC06F6573746962756C75;
        inPKT[368]      = 80'hC0706D20656C69742065;
        inPKT[369]      = 80'hC0716C656966656E6420;
        inPKT[370]      = 80'hC072756C747269636965;
        inPKT[371]      = 80'hC073732E205365642076;
        inPKT[372]      = 80'hC0746974616520646961;
        inPKT[373]      = 80'hC0756D206D6178696D75;
        inPKT[374]      = 80'hC076732C2073656D7065;
        inPKT[375]      = 80'hC07772206C6563747573;
        inPKT[376]      = 80'hC078206E65632C207661;
        inPKT[377]      = 80'hC079726975732065726F;
        inPKT[378]      = 80'hC07A732E205574206575;
        inPKT[379]      = 80'hC07B20616363756D7361;
        inPKT[380]      = 80'hC07C6E206C6967756C61;
        inPKT[381]      = 80'hC07D2E2053757370656E;
        inPKT[382]      = 80'hC07E6469737365206A75;
        inPKT[383]      = 80'hC07F73746F2072697375;
        inPKT[384]      = 80'hC080732C20736F6C6C69;
        inPKT[385]      = 80'hC0816369747564696E20;
        inPKT[386]      = 80'hC08273697420616D6574;
        inPKT[387]      = 80'hC0832068656E64726572;
        inPKT[388]      = 80'hC084697420696E2C2073;
        inPKT[389]      = 80'hC08563656C6572697371;
        inPKT[390]      = 80'hC0867565206567657420;
        inPKT[391]      = 80'hC0876D692E204E616D20;
        inPKT[392]      = 80'hC08870656C6C656E7465;
        inPKT[393]      = 80'hC0897371756520766568;
        inPKT[394]      = 80'hC08A6963756C61206469;
        inPKT[395]      = 80'hC08B676E697373696D2E;
        inPKT[396]      = 80'hC08C205365642073656D;
        inPKT[397]      = 80'hC08D7065722061756775;
        inPKT[398]      = 80'hC08E6520766974616520;
        inPKT[399]      = 80'hC08F696D706572646965;
        inPKT[400]      = 80'hC0907420736F6C6C6963;
        inPKT[401]      = 80'hC09169747564696E2E20;
        inPKT[402]      = 80'hC092566976616D757320;
        inPKT[403]      = 80'hC093616C697175616D20;
        inPKT[404]      = 80'hC0946D61676E61207669;
        inPKT[405]      = 80'hC095746165206C616375;
        inPKT[406]      = 80'hC096732072686F6E6375;
        inPKT[407]      = 80'hC0977320656C656D656E;
        inPKT[408]      = 80'hC09874756D2E20447569;
        inPKT[409]      = 80'hC099732065726F732076;
        inPKT[410]      = 80'hC09A656C69742C206C75;
        inPKT[411]      = 80'hC09B6374757320616320;
        inPKT[412]      = 80'hC09C706F72747469746F;
        inPKT[413]      = 80'hC09D72207365642C2065;
        inPKT[414]      = 80'hC09E6C656D656E74756D;
        inPKT[415]      = 80'hC09F206567657420656C;
        inPKT[416]      = 80'hC0A069742E0D0A0D0A53;
        inPKT[417]      = 80'hC0A1656420636F6E7661;
        inPKT[418]      = 80'hC0A26C6C6973206E6571;
        inPKT[419]      = 80'hC0A375652076656C2069;
        inPKT[420]      = 80'hC0A46E74657264756D20;
        inPKT[421]      = 80'hC0A56D61747469732E20;
        inPKT[422]      = 80'hC0A644756973206C616F;
        inPKT[423]      = 80'hC0A77265657420656E69;
        inPKT[424]      = 80'hC0A86D2076656C207465;
        inPKT[425]      = 80'hC0A96D706F7220626962;
        inPKT[426]      = 80'hC0AA656E64756D2E2045;
        inPKT[427]      = 80'hC0AB7469616D20736F64;
        inPKT[428]      = 80'hC0AC616C6573206D6175;
        inPKT[429]      = 80'hC0AD726973206E656320;
        inPKT[430]      = 80'hC0AE6D61676E6120626C;
        inPKT[431]      = 80'hC0AF616E6469742C2061;
        inPKT[432]      = 80'hC0B074206D6174746973;
        inPKT[433]      = 80'hC0B1206E756C6C612063;
        inPKT[434]      = 80'hC0B26F6E736571756174;
        inPKT[435]      = 80'hC0B32E20496E74657264;
        inPKT[436]      = 80'hC0B4756D206574206D61;
        inPKT[437]      = 80'hC0B56C65737561646120;
        inPKT[438]      = 80'hC0B666616D6573206163;
        inPKT[439]      = 80'hC0B720616E7465206970;
        inPKT[440]      = 80'hC0B873756D207072696D;
        inPKT[441]      = 80'hC0B9697320696E206661;
        inPKT[442]      = 80'hC0BA7563696275732E20;
        inPKT[443]      = 80'hC0BB566976616D757320;
        inPKT[444]      = 80'hC0BC6C616F7265657420;
        inPKT[445]      = 80'hC0BD756C747269636573;
        inPKT[446]      = 80'hC0BE2073656D7065722E;
        inPKT[447]      = 80'hC0BF20566976616D7573;
        inPKT[448]      = 80'hC0C0206E6F6E20647569;
        inPKT[449]      = 80'hC0C12073697420616D65;
        inPKT[450]      = 80'hC0C27420647569207375;
        inPKT[451]      = 80'hC0C37363697069742075;
        inPKT[452]      = 80'hC0C46C6C616D636F7270;
        inPKT[453]      = 80'hC0C565722E204D617572;
        inPKT[454]      = 80'hC0C66973206574206C69;
        inPKT[455]      = 80'hC0C767756C6120616C69;
        inPKT[456]      = 80'hC0C8717565742C206375;
        inPKT[457]      = 80'hC0C972737573206D6167;
        inPKT[458]      = 80'hC0CA6E612061632C2073;
        inPKT[459]      = 80'hC0CB63656C6572697371;
        inPKT[460]      = 80'hC0CC7565206A7573746F;
        inPKT[461]      = 80'hC0CD2E20416C69717561;
        inPKT[462]      = 80'hC0CE6D2076656C206469;
        inPKT[463]      = 80'hC0CF676E697373696D20;
        inPKT[464]      = 80'hC0D06469616D2E204475;
        inPKT[465]      = 80'hC0D169732076656C206E;
        inPKT[466]      = 80'hC0D2756E632065742061;
        inPKT[467]      = 80'hC0D37263752070686172;
        inPKT[468]      = 80'hC0D46574726120727574;
        inPKT[469]      = 80'hC0D572756D2071756973;
        inPKT[470]      = 80'hC0D62061742065726174;
        inPKT[471]      = 80'hC0D72E0D0A0D0A496E20;
        inPKT[472]      = 80'hC0D86F726369206C6563;
        inPKT[473]      = 80'hC0D97475732C20706F72;
        inPKT[474]      = 80'hC0DA747469746F722076;
        inPKT[475]      = 80'hC0DB656C20746F72746F;
        inPKT[476]      = 80'hC0DC72206C6F626F7274;
        inPKT[477]      = 80'hC0DD69732C2066657567;
        inPKT[478]      = 80'hC0DE6961742065676573;
        inPKT[479]      = 80'hC0DF746173206469616D;
        inPKT[480]      = 80'hC0E02E2043726173206C;
        inPKT[481]      = 80'hC0E1696265726F207075;
        inPKT[482]      = 80'hC0E27275732C206C6F62;
        inPKT[483]      = 80'hC0E36F72746973206575;
        inPKT[484]      = 80'hC0E4206E69736C206174;
        inPKT[485]      = 80'hC0E52C20616C69717565;
        inPKT[486]      = 80'hC0E67420766573746962;
        inPKT[487]      = 80'hC0E7756C756D206C6563;
        inPKT[488]      = 80'hC0E87475732E20557420;
        inPKT[489]      = 80'hC0E9696D706572646965;
        inPKT[490]      = 80'hC0EA74206469616D2073;
        inPKT[491]      = 80'hC0EB697420616D657420;
        inPKT[492]      = 80'hC0EC6E756C6C61206865;
        inPKT[493]      = 80'hC0ED6E6472657269742C;
        inPKT[494]      = 80'hC0EE2073656420766976;
        inPKT[495]      = 80'hC0EF6572726120657261;
        inPKT[496]      = 80'hC0F07420636F6E76616C;
        inPKT[497]      = 80'hC0F16C69732E20557420;
        inPKT[498]      = 80'hC0F26D6178696D75732C;
        inPKT[499]      = 80'hC0F3206C6967756C6120;
        inPKT[500]      = 80'hC0F473697420616D6574;
        inPKT[501]      = 80'hC0F52065666669636974;
        inPKT[502]      = 80'hC0F67572206D6178696D;
        inPKT[503]      = 80'hC0F775732C2073617069;
        inPKT[504]      = 80'hC0F8656E206C6F72656D;
        inPKT[505]      = 80'hC0F920636F6E67756520;
        inPKT[506]      = 80'hC0FA6F64696F2C20756C;
        inPKT[507]      = 80'hC0FB7472696365732066;
        inPKT[508]      = 80'hC0FC65726D656E74756D;
        inPKT[509]      = 80'hC0FD206E756E63206D61;
        inPKT[510]      = 80'hC0FE75726973206E6563;
        inPKT[511]      = 80'hC0FF206E6962682E2043;
        inPKT[512]      = 80'hC0007572616269747572;
        inPKT[513]      = 80'hC0012072697375732064;
        inPKT[514]      = 80'hC0026F6C6F722C20756C;
        inPKT[515]      = 80'hC0037472696369657320;
        inPKT[516]      = 80'hC0047175697320647569;
        inPKT[517]      = 80'hC0052076697461652C20;
        inPKT[518]      = 80'hC006616C697175657420;
        inPKT[519]      = 80'hC00770756C76696E6172;
        inPKT[520]      = 80'hC00820656C69742E2045;
        inPKT[521]      = 80'hC0097469616D20736167;
        inPKT[522]      = 80'hC00A6974746973206970;
        inPKT[523]      = 80'hC00B73756D206D617373;
        inPKT[524]      = 80'hC00C612C207669746165;
        inPKT[525]      = 80'hC00D20636F6E64696D65;
        inPKT[526]      = 80'hC00E6E74756D2066656C;
        inPKT[527]      = 80'hC00F697320616C697175;
        inPKT[528]      = 80'hC01065742065752E2050;
        inPKT[529]      = 80'hC01172616573656E7420;
        inPKT[530]      = 80'hC012766F6C7574706174;
        inPKT[531]      = 80'hC01320656C6974206665;
        inPKT[532]      = 80'hC0147567696174207475;
        inPKT[533]      = 80'hC015727069732074656D;
        inPKT[534]      = 80'hC016706F722068656E64;
        inPKT[535]      = 80'hC01772657269742E2041;
        inPKT[536]      = 80'hC018656E65616E206163;
        inPKT[537]      = 80'hC01963756D73616E2C20;
        inPKT[538]      = 80'hC01A65726F7320656765;
        inPKT[539]      = 80'hC01B7420696D70657264;
        inPKT[540]      = 80'hC01C6965742070656C6C;
        inPKT[541]      = 80'hC01D656E746573717565;
        inPKT[542]      = 80'hC01E2C2073656D206D69;
        inPKT[543]      = 80'hC01F2076697665727261;
        inPKT[544]      = 80'hC02020656C69742C2073;
        inPKT[545]      = 80'hC0216F64616C65732070;
        inPKT[546]      = 80'hC022756C76696E617220;
        inPKT[547]      = 80'hC0237269737573206A75;
        inPKT[548]      = 80'hC02473746F2071756973;
        inPKT[549]      = 80'hC02520616E74652E2044;
        inPKT[550]      = 80'hC0266F6E656320656C65;
        inPKT[551]      = 80'hC0276D656E74756D2065;
        inPKT[552]      = 80'hC028737420657520696D;
        inPKT[553]      = 80'hC0297065726469657420;
        inPKT[554]      = 80'hC02A756C747269636965;
        inPKT[555]      = 80'hC02B732E2050656C6C65;
        inPKT[556]      = 80'hC02C6E74657371756520;
        inPKT[557]      = 80'hC02D756C747269636573;
        inPKT[558]      = 80'hC02E206E65717565206E;
        inPKT[559]      = 80'hC02F6563206C656F206C;
        inPKT[560]      = 80'hC030616F726565742C20;
        inPKT[561]      = 80'hC031612070756C76696E;
        inPKT[562]      = 80'hC0326172206475692075;
        inPKT[563]      = 80'hC0336C6C616D636F7270;
        inPKT[564]      = 80'hC03465722E204D6F7262;
        inPKT[565]      = 80'hC0356920657569736D6F;
        inPKT[566]      = 80'hC036642C206D65747573;
        inPKT[567]      = 80'hC03720696420616C6971;
        inPKT[568]      = 80'hC03875657420616C6971;
        inPKT[569]      = 80'hC03975616D2C206C6F72;
        inPKT[570]      = 80'hC03A656D206A7573746F;
        inPKT[571]      = 80'hC03B20666163696C6973;
        inPKT[572]      = 80'hC03C697320646F6C6F72;
        inPKT[573]      = 80'hC03D2C206E6F6E206461;
        inPKT[574]      = 80'hC03E7069627573206572;
        inPKT[575]      = 80'hC03F6174206D69207669;
        inPKT[576]      = 80'hC040746165206E756E63;
        inPKT[577]      = 80'hC0412E20536564206574;
        inPKT[578]      = 80'hC0422065726F73206120;
        inPKT[579]      = 80'hC04373617069656E2061;
        inPKT[580]      = 80'hC0447563746F7220756C;
        inPKT[581]      = 80'hC0457472696365732E20;
        inPKT[582]      = 80'hC0465175697371756520;
        inPKT[583]      = 80'hC0477175697320636F6E;
        inPKT[584]      = 80'hC04864696D656E74756D;
        inPKT[585]      = 80'hC049206A7573746F2E20;
        inPKT[586]      = 80'hC04A446F6E6563207465;
        inPKT[587]      = 80'hC04B6C6C7573206A7573;
        inPKT[588]      = 80'hC04C746F2C20706F7274;
        inPKT[589]      = 80'hC04D6120717569732073;
        inPKT[590]      = 80'hC04E617069656E20612C;
        inPKT[591]      = 80'hC04F20696D7065726469;
        inPKT[592]      = 80'hC0506574206C75637475;
        inPKT[593]      = 80'hC05173206573742E204D;
        inPKT[594]      = 80'hC0526F72626920626962;
        inPKT[595]      = 80'hC053656E64756D206E69;
        inPKT[596]      = 80'hC054736C20616E74652C;
        inPKT[597]      = 80'hC0552065752064696374;
        inPKT[598]      = 80'hC056756D206E65717565;
        inPKT[599]      = 80'hC05720696D7065726469;
        inPKT[600]      = 80'hC05865742065742E2050;
        inPKT[601]      = 80'hC059686173656C6C7573;
        inPKT[602]      = 80'hC05A2071756973207361;
        inPKT[603]      = 80'hC05B7069656E20617567;
        inPKT[604]      = 80'hC05C75652E0D0A0D0A49;
        inPKT[605]      = 80'hC05D6E74656765722069;
        inPKT[606]      = 80'hC05E6E2073617069656E;
        inPKT[607]      = 80'hC05F20746F72746F722E;
        inPKT[608]      = 80'hC060204D617572697320;
        inPKT[609]      = 80'hC061657520656E696D20;
        inPKT[610]      = 80'hC0626D692E2056697661;
        inPKT[611]      = 80'hC0636D7573206C616369;
        inPKT[612]      = 80'hC0646E6961206D61676E;
        inPKT[613]      = 80'hC06561206E6563206573;
        inPKT[614]      = 80'hC0667420656C65696665;
        inPKT[615]      = 80'hC0676E642C2061742063;
        inPKT[616]      = 80'hC0686F6E67756520616E;
        inPKT[617]      = 80'hC069746520706C616365;
        inPKT[618]      = 80'hC06A7261742E20437261;
        inPKT[619]      = 80'hC06B7320736564206665;
        inPKT[620]      = 80'hC06C726D656E74756D20;
        inPKT[621]      = 80'hC06D76656C69742E2053;
        inPKT[622]      = 80'hC06E6564206C616F7265;
        inPKT[623]      = 80'hC06F6574206C69626572;
        inPKT[624]      = 80'hC0706F20616320746F72;
        inPKT[625]      = 80'hC071746F722065756973;
        inPKT[626]      = 80'hC0726D6F642C20656765;
        inPKT[627]      = 80'hC0737420766976657272;
        inPKT[628]      = 80'hC0746120656C69742064;
        inPKT[629]      = 80'hC075696374756D2E2053;
        inPKT[630]      = 80'hC076757370656E646973;
        inPKT[631]      = 80'hC077736520756C747269;
        inPKT[632]      = 80'hC0786365732069642064;
        inPKT[633]      = 80'hC07969616D2065676574;
        inPKT[634]      = 80'hC07A20756C6C616D636F;
        inPKT[635]      = 80'hC07B727065722E205072;
        inPKT[636]      = 80'hC07C616573656E74206D;
        inPKT[637]      = 80'hC07D6F6C6C6973207465;
        inPKT[638]      = 80'hC07E6D70757320746F72;
        inPKT[639]      = 80'hC07F746F722069642063;
        inPKT[640]      = 80'hC0806F6E736571756174;
        inPKT[641]      = 80'hC0812E204E616D206F72;
        inPKT[642]      = 80'hC0826E61726520616320;
        inPKT[643]      = 80'hC0836E65717565207175;
        inPKT[644]      = 80'hC084697320756C747269;
        inPKT[645]      = 80'hC0856365732E20447569;
        inPKT[646]      = 80'hC086732061742076656E;
        inPKT[647]      = 80'hC087656E617469732064;
        inPKT[648]      = 80'hC08869616D2C206D6F6C;
        inPKT[649]      = 80'hC089657374696520636F;
        inPKT[650]      = 80'hC08A6E73657175617420;
        inPKT[651]      = 80'hC08B6E756E632E204D61;
        inPKT[652]      = 80'hC08C6563656E6173206E;
        inPKT[653]      = 80'hC08D6563206C61637573;
        inPKT[654]      = 80'hC08E2076656C69742E20;
        inPKT[655]      = 80'hC08F5175697371756520;
        inPKT[656]      = 80'hC0906772617669646120;
        inPKT[657]      = 80'hC0916469616D206E6563;
        inPKT[658]      = 80'hC0922073656D20737573;
        inPKT[659]      = 80'hC09363697069742C2073;
        inPKT[660]      = 80'hC0946564206C6163696E;
        inPKT[661]      = 80'hC0956961207175616D20;
        inPKT[662]      = 80'hC09670756C76696E6172;
        inPKT[663]      = 80'hC0972E0D0A0D0A496E20;
        inPKT[664]      = 80'hC098696D706572646965;
        inPKT[665]      = 80'hC099742065726F73206F;
        inPKT[666]      = 80'hC09A726E617265206578;
        inPKT[667]      = 80'hC09B207665686963756C;
        inPKT[668]      = 80'hC09C612C20657420696E;
        inPKT[669]      = 80'hC09D74657264756D206C;
        inPKT[670]      = 80'hC09E6163757320637572;
        inPKT[671]      = 80'hC09F7375732E204D6175;
        inPKT[672]      = 80'hC0A07269732065742073;
        inPKT[673]      = 80'hC0A1656D706572206175;
        inPKT[674]      = 80'hC0A26775652C20766974;
        inPKT[675]      = 80'hC0A36165206D6F6C6C69;
        inPKT[676]      = 80'hC0A473206C6563747573;
        inPKT[677]      = 80'hC0A52E20517569737175;
        inPKT[678]      = 80'hC0A6652073697420616D;
        inPKT[679]      = 80'hC0A76574206C656F2071;
        inPKT[680]      = 80'hC0A875697320616E7465;
        inPKT[681]      = 80'hC0A92063757273757320;
        inPKT[682]      = 80'hC0AA616C69717565742E;
        inPKT[683]      = 80'hC0AB204D617572697320;
        inPKT[684]      = 80'hC0AC7068617265747261;
        inPKT[685]      = 80'hC0AD2076656C69742076;
        inPKT[686]      = 80'hC0AE656C20626962656E;
        inPKT[687]      = 80'hC0AF64756D2074656D70;
        inPKT[688]      = 80'hC0B075732E20496E2068;
        inPKT[689]      = 80'hC0B16163206861626974;
        inPKT[690]      = 80'hC0B26173736520706C61;
        inPKT[691]      = 80'hC0B37465612064696374;
        inPKT[692]      = 80'hC0B4756D73742E20496E;
        inPKT[693]      = 80'hC0B52076657374696275;
        inPKT[694]      = 80'hC0B66C756D2C2075726E;
        inPKT[695]      = 80'hC0B76120657420736F6C;
        inPKT[696]      = 80'hC0B86C69636974756469;
        inPKT[697]      = 80'hC0B96E2070756C76696E;
        inPKT[698]      = 80'hC0BA61722C206E69736C;
        inPKT[699]      = 80'hC0BB2065737420656666;
        inPKT[700]      = 80'hC0BC6963697475722071;
        inPKT[701]      = 80'hC0BD75616D2C206D6F6C;
        inPKT[702]      = 80'hC0BE6C6973206C616F72;
        inPKT[703]      = 80'hC0BF6565742065726174;
        inPKT[704]      = 80'hC0C0206D692061206C6F;
        inPKT[705]      = 80'hC0C172656D2E20457469;
        inPKT[706]      = 80'hC0C2616D207574206C65;
        inPKT[707]      = 80'hC0C36F2065782E204165;
        inPKT[708]      = 80'hC0C46E65616E206D6574;
        inPKT[709]      = 80'hC0C5757320617263752C;
        inPKT[710]      = 80'hC0C620696D7065726469;
        inPKT[711]      = 80'hC0C76574206574207361;
        inPKT[712]      = 80'hC0C87069656E20696E2C;
        inPKT[713]      = 80'hC0C920617563746F7220;
        inPKT[714]      = 80'hC0CA616363756D73616E;
        inPKT[715]      = 80'hC0CB2065782E20566976;
        inPKT[716]      = 80'hC0CC616D757320706F73;
        inPKT[717]      = 80'hC0CD756572652075726E;
        inPKT[718]      = 80'hC0CE6120696420657261;
        inPKT[719]      = 80'hC0CF742072686F6E6375;
        inPKT[720]      = 80'hC0D07320666575676961;
        inPKT[721]      = 80'hC0D1742E205068617365;
        inPKT[722]      = 80'hC0D26C6C7573206D6175;
        inPKT[723]      = 80'hC0D372697320656C6974;
        inPKT[724]      = 80'hC0D42C20677261766964;
        inPKT[725]      = 80'hC0D561206575206D6F6C;
        inPKT[726]      = 80'hC0D66C6973207365642C;
        inPKT[727]      = 80'hC0D7206C616F72656574;
        inPKT[728]      = 80'hC0D82071756973206E75;
        inPKT[729]      = 80'hC0D96E632E20496E7465;
        inPKT[730]      = 80'hC0DA6765722069616375;
        inPKT[731]      = 80'hC0DB6C697320656E696D;
        inPKT[732]      = 80'hC0DC20617263752C2065;
        inPKT[733]      = 80'hC0DD676574206D617869;
        inPKT[734]      = 80'hC0DE6D7573206C656374;
        inPKT[735]      = 80'hC0DF757320766F6C7574;
        inPKT[736]      = 80'hC0E0706174206E6F6E2E;
        inPKT[737]      = 80'hC0E120496E7465726475;
        inPKT[738]      = 80'hC0E26D206574206D616C;
        inPKT[739]      = 80'hC0E36573756164612066;
        inPKT[740]      = 80'hC0E4616D657320616320;
        inPKT[741]      = 80'hC0E5616E746520697073;
        inPKT[742]      = 80'hC0E6756D207072696D69;
        inPKT[743]      = 80'hC0E77320696E20666175;
        inPKT[744]      = 80'hC0E863696275732E2044;
        inPKT[745]      = 80'hC0E96F6E656320696E20;
        inPKT[746]      = 80'hC0EA7475727069732063;
        inPKT[747]      = 80'hC0EB7572737573207475;
        inPKT[748]      = 80'hC0EC72706973206D6F6C;
        inPKT[749]      = 80'hC0ED657374696520636F;
        inPKT[750]      = 80'hC0EE6E73657175617420;
        inPKT[751]      = 80'hC0EF6174206174207269;
        inPKT[752]      = 80'hC0F07375732E0D0A0D0A;
        inPKT[753]      = 80'hC0F1446F6E6563207365;
        inPKT[754]      = 80'hC0F26D206E756E632C20;
        inPKT[755]      = 80'hC0F3636F6E7365637465;
        inPKT[756]      = 80'hC0F47475722061207465;
        inPKT[757]      = 80'hC0F56C6C757320612C20;
        inPKT[758]      = 80'hC0F6616363756D73616E;
        inPKT[759]      = 80'hC0F72070656C6C656E74;
        inPKT[760]      = 80'hC0F86573717565207075;
        inPKT[761]      = 80'hC0F97275732E20507261;
        inPKT[762]      = 80'hC0FA6573656E74206375;
        inPKT[763]      = 80'hC0FB727375732074656D;
        inPKT[764]      = 80'hC0FC706F722064617069;
        inPKT[765]      = 80'hC0FD6275732E20457469;
        inPKT[766]      = 80'hC0FE616D2076656C6974;
        inPKT[767]      = 80'hC0FF206475692C207375;
        inPKT[768]      = 80'hC0007363697069742076;
        inPKT[769]      = 80'hC0016974616520756C6C;
        inPKT[770]      = 80'hC002616D636F72706572;
        inPKT[771]      = 80'hC00320636F6D6D6F646F;
        inPKT[772]      = 80'hC0042C206C7563747573;
        inPKT[773]      = 80'hC005206469676E697373;
        inPKT[774]      = 80'hC006696D207075727573;
        inPKT[775]      = 80'hC0072E2053757370656E;
        inPKT[776]      = 80'hC008646973736520706F;
        inPKT[777]      = 80'hC00974656E74692E2049;
        inPKT[778]      = 80'hC00A6E20637572737573;
        inPKT[779]      = 80'hC00B20697073756D2074;
        inPKT[780]      = 80'hC00C656D706F72207175;
        inPKT[781]      = 80'hC00D616D2074696E6369;
        inPKT[782]      = 80'hC00E64756E7420747269;
        inPKT[783]      = 80'hC00F7374697175652065;
        inPKT[784]      = 80'hC0106765742073656420;
        inPKT[785]      = 80'hC0116D692E2045746961;
        inPKT[786]      = 80'hC0126D2074696E636964;
        inPKT[787]      = 80'hC013756E74207175616D;
        inPKT[788]      = 80'hC0142075742076656C69;
        inPKT[789]      = 80'hC0157420747269737469;
        inPKT[790]      = 80'hC016717565206C6F626F;
        inPKT[791]      = 80'hC017727469732E20446F;
        inPKT[792]      = 80'hC0186E6563206E657175;
        inPKT[793]      = 80'hC01965206D692C20736F;
        inPKT[794]      = 80'hC01A6C6C696369747564;
        inPKT[795]      = 80'hC01B696E207369742061;
        inPKT[796]      = 80'hC01C6D657420656E696D;
        inPKT[797]      = 80'hC01D20696E2C20656666;
        inPKT[798]      = 80'hC01E6963697475722070;
        inPKT[799]      = 80'hC01F6F7274612073656D;
        inPKT[800]      = 80'hC0202E20437572616269;
        inPKT[801]      = 80'hC0217475722061742070;
        inPKT[802]      = 80'hC022756C76696E617220;
        inPKT[803]      = 80'hC0236E6962682E205065;
        inPKT[804]      = 80'hC0246C6C656E74657371;
        inPKT[805]      = 80'hC02575652076656C2061;
        inPKT[806]      = 80'hC0266C697175616D206A;
        inPKT[807]      = 80'hC0277573746F2E20416C;
        inPKT[808]      = 80'hC028697175616D206572;
        inPKT[809]      = 80'hC029617420766F6C7574;
        inPKT[810]      = 80'hC02A7061742E20536564;
        inPKT[811]      = 80'hC02B207365642076656C;
        inPKT[812]      = 80'hC02C6974206E6973692E;
        inPKT[813]      = 80'hC02D2046757363652063;
        inPKT[814]      = 80'hC02E757273757320696E;
        inPKT[815]      = 80'hC02F74657264756D206C;
        inPKT[816]      = 80'hC0306F626F727469732E;
        inPKT[817]      = 80'hC0310D0A0D0A50726165;
        inPKT[818]      = 80'hC03273656E7420706F73;
        inPKT[819]      = 80'hC0337565726520696E20;
        inPKT[820]      = 80'hC0346572617420736564;
        inPKT[821]      = 80'hC0352072686F6E637573;
        inPKT[822]      = 80'hC0362E20446F6E656320;
        inPKT[823]      = 80'hC0376575206573742065;
        inPKT[824]      = 80'hC03874206C6563747573;
        inPKT[825]      = 80'hC039206C6163696E6961;
        inPKT[826]      = 80'hC03A2070756C76696E61;
        inPKT[827]      = 80'hC03B722E204675736365;
        inPKT[828]      = 80'hC03C2076656E656E6174;
        inPKT[829]      = 80'hC03D6973206572617420;
        inPKT[830]      = 80'hC03E75726E612C206574;
        inPKT[831]      = 80'hC03F2073616769747469;
        inPKT[832]      = 80'hC040732073617069656E;
        inPKT[833]      = 80'hC0412076617269757320;
        inPKT[834]      = 80'hC04273697420616D6574;
        inPKT[835]      = 80'hC0432E20467573636520;
        inPKT[836]      = 80'hC0446475692065726174;
        inPKT[837]      = 80'hC0452C20766976657272;
        inPKT[838]      = 80'hC04661207574206C6F62;
        inPKT[839]      = 80'hC0476F72746973207365;
        inPKT[840]      = 80'hC048642C20666163696C;
        inPKT[841]      = 80'hC0496973697320717569;
        inPKT[842]      = 80'hC04A73206D657475732E;
        inPKT[843]      = 80'hC04B204D6F7262692067;
        inPKT[844]      = 80'hC04C726176696461206D;
        inPKT[845]      = 80'hC04D61737361206E6F6E;
        inPKT[846]      = 80'hC04E207072657469756D;
        inPKT[847]      = 80'hC04F2066696E69627573;
        inPKT[848]      = 80'hC0502E204D616563656E;
        inPKT[849]      = 80'hC0516173206C6F72656D;
        inPKT[850]      = 80'hC052207475727069732C;
        inPKT[851]      = 80'hC0532063757273757320;
        inPKT[852]      = 80'hC05475742076656C6974;
        inPKT[853]      = 80'hC05520612C2061636375;
        inPKT[854]      = 80'hC0566D73616E2074696E;
        inPKT[855]      = 80'hC057636964756E74206F;
        inPKT[856]      = 80'hC05864696F2E2050726F;
        inPKT[857]      = 80'hC059696E20656C697420;
        inPKT[858]      = 80'hC05A76656C69742C2065;
        inPKT[859]      = 80'hC05B6C656D656E74756D;
        inPKT[860]      = 80'hC05C2076656C20696163;
        inPKT[861]      = 80'hC05D756C69732065752C;
        inPKT[862]      = 80'hC05E20636F6E64696D65;
        inPKT[863]      = 80'hC05F6E74756D20657420;
        inPKT[864]      = 80'hC06075726E612E205665;
        inPKT[865]      = 80'hC06173746962756C756D;
        inPKT[866]      = 80'hC062206E656320657820;
        inPKT[867]      = 80'hC0636F7263692E204675;
        inPKT[868]      = 80'hC064736365206174206C;
        inPKT[869]      = 80'hC0656F72656D20617420;
        inPKT[870]      = 80'hC0666C6163757320696E;
        inPKT[871]      = 80'hC06774657264756D2064;
        inPKT[872]      = 80'hC068696374756D2E2041;
        inPKT[873]      = 80'hC0696C697175616D2073;
        inPKT[874]      = 80'hC06A656D70657220766F;
        inPKT[875]      = 80'hC06B6C75747061742070;
        inPKT[876]      = 80'hC06C6F73756572652E20;
        inPKT[877]      = 80'hC06D4E756C6C616D2076;
        inPKT[878]      = 80'hC06E656C20647569206C;
        inPKT[879]      = 80'hC06F6163696E69612C20;
        inPKT[880]      = 80'hC07070656C6C656E7465;
        inPKT[881]      = 80'hC0717371756520657820;
        inPKT[882]      = 80'hC072717569732C20756C;
        inPKT[883]      = 80'hC0736C616D636F727065;
        inPKT[884]      = 80'hC07472206F7263692E20;
        inPKT[885]      = 80'hC0754372617320666572;
        inPKT[886]      = 80'hC0766D656E74756D2C20;
        inPKT[887]      = 80'hC0776C61637573207574;
        inPKT[888]      = 80'hC0782070756C76696E61;
        inPKT[889]      = 80'hC0797220636F6E736571;
        inPKT[890]      = 80'hC07A7561742C206D6574;
        inPKT[891]      = 80'hC07B7573207361706965;
        inPKT[892]      = 80'hC07C6E20656666696369;
        inPKT[893]      = 80'hC07D747572206E69736C;
        inPKT[894]      = 80'hC07E2C20696E206D6F6C;
        inPKT[895]      = 80'hC07F6573746965206E69;
        inPKT[896]      = 80'hC0807369206C69626572;
        inPKT[897]      = 80'hC0816F20696E2076656C;
        inPKT[898]      = 80'hC08269742E204D616563;
        inPKT[899]      = 80'hC083656E6173206D6173;
        inPKT[900]      = 80'hC084736120746F72746F;
        inPKT[901]      = 80'hC085722C207275747275;
        inPKT[902]      = 80'hC0866D2076656C206669;
        inPKT[903]      = 80'hC0876E69627573206174;
        inPKT[904]      = 80'hC0882C207363656C6572;
        inPKT[905]      = 80'hC0896973717565206574;
        inPKT[906]      = 80'hC08A206475692E20496E;
        inPKT[907]      = 80'hC08B206D616C65737561;
        inPKT[908]      = 80'hC08C64612C2066656C69;
        inPKT[909]      = 80'hC08D73206E6F6E206D6F;
        inPKT[910]      = 80'hC08E6C65737469652075;
        inPKT[911]      = 80'hC08F6C7472696365732C;
        inPKT[912]      = 80'hC090206C61637573206E;
        inPKT[913]      = 80'hC0916571756520657569;
        inPKT[914]      = 80'hC092736D6F642076656C;
        inPKT[915]      = 80'hC09369742C2076656C20;
        inPKT[916]      = 80'hC094696E74657264756D;
        inPKT[917]      = 80'hC095206D61676E612061;
        inPKT[918]      = 80'hC0966E74652061632065;
        inPKT[919]      = 80'hC09773742E0D0A0D0A49;
        inPKT[920]      = 80'hC0986E7465676572206F;
        inPKT[921]      = 80'hC099726E61726520696E;
        inPKT[922]      = 80'hC09A2075726E61206120;
        inPKT[923]      = 80'hC09B626962656E64756D;
        inPKT[924]      = 80'hC09C2E204E756C6C616D;
        inPKT[925]      = 80'hC09D207269737573206C;
        inPKT[926]      = 80'hC09E696265726F2C2076;
        inPKT[927]      = 80'hC09F756C707574617465;
        inPKT[928]      = 80'hC0A02076656C206D6920;
        inPKT[929]      = 80'hC0A16E65632C20626C61;
        inPKT[930]      = 80'hC0A26E64697420666575;
        inPKT[931]      = 80'hC0A36769617420746F72;
        inPKT[932]      = 80'hC0A4746F722E20496E20;
        inPKT[933]      = 80'hC0A56861632068616269;
        inPKT[934]      = 80'hC0A6746173736520706C;
        inPKT[935]      = 80'hC0A76174656120646963;
        inPKT[936]      = 80'hC0A874756D73742E2053;
        inPKT[937]      = 80'hC0A9757370656E646973;
        inPKT[938]      = 80'hC0AA7365207669746165;
        inPKT[939]      = 80'hC0AB20657374206A7573;
        inPKT[940]      = 80'hC0AC746F2E204E756E63;
        inPKT[941]      = 80'hC0AD20696420646F6C6F;
        inPKT[942]      = 80'hC0AE7220646170696275;
        inPKT[943]      = 80'hC0AF732C207661726975;
        inPKT[944]      = 80'hC0B07320726973757320;
        inPKT[945]      = 80'hC0B176697461652C2066;
        inPKT[946]      = 80'hC0B26163696C69736973;
        inPKT[947]      = 80'hC0B3206E6973692E2051;
        inPKT[948]      = 80'hC0B4756973717565206E;
        inPKT[949]      = 80'hC0B56973692065782C20;
        inPKT[950]      = 80'hC0B676756C7075746174;
        inPKT[951]      = 80'hC0B76520736564207363;
        inPKT[952]      = 80'hC0B8656C657269737175;
        inPKT[953]      = 80'hC0B9652076656C2C2070;
        inPKT[954]      = 80'hC0BA72657469756D2061;
        inPKT[955]      = 80'hC0BB74207175616D2E20;
        inPKT[956]      = 80'hC0BC4372617320736365;
        inPKT[957]      = 80'hC0BD6C65726973717565;
        inPKT[958]      = 80'hC0BE206120616E746520;
        inPKT[959]      = 80'hC0BF616320736F6C6C69;
        inPKT[960]      = 80'hC0C06369747564696E2E;
        inPKT[961]      = 80'hC0C10D0A0D0A41656E65;
        inPKT[962]      = 80'hC0C2616E207072657469;
        inPKT[963]      = 80'hC0C3756D2C206C6F7265;
        inPKT[964]      = 80'hC0C46D20736564206661;
        inPKT[965]      = 80'hC0C563696C6973697320;
        inPKT[966]      = 80'hC0C676656E656E617469;
        inPKT[967]      = 80'hC0C7732C206D69206E75;
        inPKT[968]      = 80'hC0C86E632076756C7075;
        inPKT[969]      = 80'hC0C97461746520616E74;
        inPKT[970]      = 80'hC0CA652C207365642070;
        inPKT[971]      = 80'hC0CB656C6C656E746573;
        inPKT[972]      = 80'hC0CC7175652066656C69;
        inPKT[973]      = 80'hC0CD732065726F732073;
        inPKT[974]      = 80'hC0CE6564206E756E632E;
        inPKT[975]      = 80'hC0CF2056657374696275;
        inPKT[976]      = 80'hC0D06C756D20616E7465;
        inPKT[977]      = 80'hC0D120697073756D2070;
        inPKT[978]      = 80'hC0D272696D697320696E;
        inPKT[979]      = 80'hC0D32066617563696275;
        inPKT[980]      = 80'hC0D473206F726369206C;
        inPKT[981]      = 80'hC0D57563747573206574;
        inPKT[982]      = 80'hC0D620756C7472696365;
        inPKT[983]      = 80'hC0D77320706F73756572;
        inPKT[984]      = 80'hC0D86520637562696C69;
        inPKT[985]      = 80'hC0D9612043757261653B;
        inPKT[986]      = 80'hC0DA2050686173656C6C;
        inPKT[987]      = 80'hC0DB757320636F6E7365;
        inPKT[988]      = 80'hC0DC717561742076756C;
        inPKT[989]      = 80'hC0DD707574617465206F;
        inPKT[990]      = 80'hC0DE7263692076656C20;
        inPKT[991]      = 80'hC0DF766F6C7574706174;
        inPKT[992]      = 80'hC0E02E20416C69717561;
        inPKT[993]      = 80'hC0E16D20657261742076;
        inPKT[994]      = 80'hC0E26F6C75747061742E;
        inPKT[995]      = 80'hC0E320446F6E65632066;
        inPKT[996]      = 80'hC0E46163696C69736973;
        inPKT[997]      = 80'hC0E52C206D61676E6120;
        inPKT[998]      = 80'hC0E661742074696E6369;
        inPKT[999]      = 80'hC0E764756E74206D6F6C;
        inPKT[1000]     = 80'hC0E86C69732C206D6920;
        inPKT[1001]     = 80'hC0E966656C6973207075;
        inPKT[1002]     = 80'hC0EA6C76696E61722065;
        inPKT[1003]     = 80'hC0EB6C69742C20617420;
        inPKT[1004]     = 80'hC0EC73656D7065722074;
        inPKT[1005]     = 80'hC0ED656C6C7573206578;
        inPKT[1006]     = 80'hC0EE20736F6C6C696369;
        inPKT[1007]     = 80'hC0EF747564696E20646F;
        inPKT[1008]     = 80'hC0F06C6F722E20517569;
        inPKT[1009]     = 80'hC0F17371756520636F6E;
        inPKT[1010]     = 80'hC0F264696D656E74756D;
        inPKT[1011]     = 80'hC0F32073617069656E20;
        inPKT[1012]     = 80'hC0F473656420706C6163;
        inPKT[1013]     = 80'hC0F56572617420706C61;
        inPKT[1014]     = 80'hC0F663657261742E2050;
        inPKT[1015]     = 80'hC0F7656C6C656E746573;
        inPKT[1016]     = 80'hC0F871756520696D7065;
        inPKT[1017]     = 80'hC0F97264696574206172;
        inPKT[1018]     = 80'hC0FA6375206573742C20;
        inPKT[1019]     = 80'hC0FB6567657420736F6C;
        inPKT[1020]     = 80'hC0FC6C69636974756469;
        inPKT[1021]     = 80'hC0FD6E2073656D206469;
        inPKT[1022]     = 80'hC0FE6374756D2061742E;
        inPKT[1023]     = 80'hC0FF2053656420736564;
        inPKT[1024]     = 80'hC000206E697369206E65;
        inPKT[1025]     = 80'hC0017175652E20537573;
        inPKT[1026]     = 80'hC00270656E6469737365;
        inPKT[1027]     = 80'hC003206D616C65737561;
        inPKT[1028]     = 80'hC0046461206D65747573;
        inPKT[1029]     = 80'hC005206E6F6E20746F72;
        inPKT[1030]     = 80'hC006746F7220636F6E67;
        inPKT[1031]     = 80'hC007756520756C6C616D;
        inPKT[1032]     = 80'hC008636F727065722E20;
        inPKT[1033]     = 80'hC009566976616D757320;
        inPKT[1034]     = 80'hC00A70656C6C656E7465;
        inPKT[1035]     = 80'hC00B7371756520717561;
        inPKT[1036]     = 80'hC00C6D207574206D6173;
        inPKT[1037]     = 80'hC00D736120626962656E;
        inPKT[1038]     = 80'hC00E64756D2064696374;
        inPKT[1039]     = 80'hC00F756D2E20496E2063;
        inPKT[1040]     = 80'hC0107572737573206174;
        inPKT[1041]     = 80'hC011206D617373612076;
        inPKT[1042]     = 80'hC0126974616520736365;
        inPKT[1043]     = 80'hC0136C65726973717565;
        inPKT[1044]     = 80'hC0142E204D616563656E;
        inPKT[1045]     = 80'hC0156173206964207465;
        inPKT[1046]     = 80'hC0166D707573206E6962;
        inPKT[1047]     = 80'hC017682E20496E206D69;
        inPKT[1048]     = 80'hC0182076656C69742C20;
        inPKT[1049]     = 80'hC019636F6E6775652061;
        inPKT[1050]     = 80'hC01A2066696E69627573;
        inPKT[1051]     = 80'hC01B2061742C206D616C;
        inPKT[1052]     = 80'hC01C657375616461206E;
        inPKT[1053]     = 80'hC01D65632073656D2E20;
        inPKT[1054]     = 80'hC01E50656C6C656E7465;
        inPKT[1055]     = 80'hC01F73717565206C6163;
        inPKT[1056]     = 80'hC020696E696120636F6E;
        inPKT[1057]     = 80'hC02164696D656E74756D;
        inPKT[1058]     = 80'hC0222076756C70757461;
        inPKT[1059]     = 80'hC02374652E2056697661;
        inPKT[1060]     = 80'hC0246D7573206E6F6E20;
        inPKT[1061]     = 80'hC0256E69626820696420;
        inPKT[1062]     = 80'hC02673656D2074656D70;
        inPKT[1063]     = 80'hC027757320696163756C;
        inPKT[1064]     = 80'hC02869732E2051756973;
        inPKT[1065]     = 80'hC0297175652076617269;
        inPKT[1066]     = 80'hC02A7573206E69626820;
        inPKT[1067]     = 80'hC02B76656C2070757275;
        inPKT[1068]     = 80'hC02C732064696374756D;
        inPKT[1069]     = 80'hC02D2074656D706F7220;
        inPKT[1070]     = 80'hC02E76656C2065752061;
        inPKT[1071]     = 80'hC02F7263752E0D0A0D0A;
        inPKT[1072]     = 80'hC03050686173656C6C75;
        inPKT[1073]     = 80'hC031732072757472756D;
        inPKT[1074]     = 80'hC032206C6967756C6120;
        inPKT[1075]     = 80'hC0336E756E632C206174;
        inPKT[1076]     = 80'hC0342066657567696174;
        inPKT[1077]     = 80'hC0352072697375732066;
        inPKT[1078]     = 80'hC03672696E67696C6C61;
        inPKT[1079]     = 80'hC0372076656C2E204372;
        inPKT[1080]     = 80'hC0386173207361706965;
        inPKT[1081]     = 80'hC0396E206D6175726973;
        inPKT[1082]     = 80'hC03A2C20766568696375;
        inPKT[1083]     = 80'hC03B6C61207574207268;
        inPKT[1084]     = 80'hC03C6F6E637573206575;
        inPKT[1085]     = 80'hC03D69736D6F642C206D;
        inPKT[1086]     = 80'hC03E616C657375616461;
        inPKT[1087]     = 80'hC03F206E6F6E20717561;
        inPKT[1088]     = 80'hC0406D2E205365642064;
        inPKT[1089]     = 80'hC04169676E697373696D;
        inPKT[1090]     = 80'hC042206F726E61726520;
        inPKT[1091]     = 80'hC0436D6178696D75732E;
        inPKT[1092]     = 80'hC0442043757261626974;
        inPKT[1093]     = 80'hC0457572207175697320;
        inPKT[1094]     = 80'hC0466C6967756C61206C;
        inPKT[1095]     = 80'hC047696265726F2E204C;
        inPKT[1096]     = 80'hC0486F72656D20697073;
        inPKT[1097]     = 80'hC049756D20646F6C6F72;
        inPKT[1098]     = 80'hC04A2073697420616D65;
        inPKT[1099]     = 80'hC04B742C20636F6E7365;
        inPKT[1100]     = 80'hC04C6374657475722061;
        inPKT[1101]     = 80'hC04D646970697363696E;
        inPKT[1102]     = 80'hC04E6720656C69742E20;
        inPKT[1103]     = 80'hC04F457469616D206D61;
        inPKT[1104]     = 80'hC05078696D7573206665;
        inPKT[1105]     = 80'hC0516C69732073656420;
        inPKT[1106]     = 80'hC05264756920706C6163;
        inPKT[1107]     = 80'hC0536572617420706F72;
        inPKT[1108]     = 80'hC05474612E204D6F7262;
        inPKT[1109]     = 80'hC055692073656420626C;
        inPKT[1110]     = 80'hC056616E646974206C65;
        inPKT[1111]     = 80'hC057637475732C206120;
        inPKT[1112]     = 80'hC058756C6C616D636F72;
        inPKT[1113]     = 80'hC059706572206E657175;
        inPKT[1114]     = 80'hC05A652E205365642069;
        inPKT[1115]     = 80'hC05B6E206E697369206D;
        inPKT[1116]     = 80'hC05C617373612E20446F;
        inPKT[1117]     = 80'hC05D6E6563206163206C;
        inPKT[1118]     = 80'hC05E7563747573206F72;
        inPKT[1119]     = 80'hC05F63692C2065752062;
        inPKT[1120]     = 80'hC0606962656E64756D20;
        inPKT[1121]     = 80'hC061646F6C6F722E2053;
        inPKT[1122]     = 80'hC0626564206D6F6C6573;
        inPKT[1123]     = 80'hC06374696520616C6971;
        inPKT[1124]     = 80'hC06475616D206E697369;
        inPKT[1125]     = 80'hC0652076656C20636F6E;
        inPKT[1126]     = 80'hC06676616C6C69732E0D;
        inPKT[1127]     = 80'hC0670A0D0A416C697175;
        inPKT[1128]     = 80'hC068616D206567657420;
        inPKT[1129]     = 80'hC069636F6E7365717561;
        inPKT[1130]     = 80'hC06A74206C616375732C;
        inPKT[1131]     = 80'hC06B207365642076656E;
        inPKT[1132]     = 80'hC06C656E61746973206C;
        inPKT[1133]     = 80'hC06D65637475732E2043;
        inPKT[1134]     = 80'hC06E7261732076656869;
        inPKT[1135]     = 80'hC06F63756C61206E6571;
        inPKT[1136]     = 80'hC070756520696E206572;
        inPKT[1137]     = 80'hC0716F73207363656C65;
        inPKT[1138]     = 80'hC072726973717565206D;
        inPKT[1139]     = 80'hC0736F6C6C69732E2050;
        inPKT[1140]     = 80'hC074656C6C656E746573;
        inPKT[1141]     = 80'hC075717565206D69206D;
        inPKT[1142]     = 80'hC07661676E612C206D6F;
        inPKT[1143]     = 80'hC0776C6573746965206E;
        inPKT[1144]     = 80'hC0786F6E20636F6E6469;
        inPKT[1145]     = 80'hC0796D656E74756D2073;
        inPKT[1146]     = 80'hC07A697420616D65742C;
        inPKT[1147]     = 80'hC07B20706F7274612076;
        inPKT[1148]     = 80'hC07C656C2075726E612E;
        inPKT[1149]     = 80'hC07D2041656E65616E20;
        inPKT[1150]     = 80'hC07E66656C6973206E75;
        inPKT[1151]     = 80'hC07F6E632C20636F6E64;
        inPKT[1152]     = 80'hC080696D656E74756D20;
        inPKT[1153]     = 80'hC081657420746F72746F;
        inPKT[1154]     = 80'hC082722074696E636964;
        inPKT[1155]     = 80'hC083756E742C20707265;
        inPKT[1156]     = 80'hC0847469756D20766172;
        inPKT[1157]     = 80'hC085697573206E756C6C;
        inPKT[1158]     = 80'hC086612E204E756E6320;
        inPKT[1159]     = 80'hC08776656C206E657175;
        inPKT[1160]     = 80'hC08865206174206C6967;
        inPKT[1161]     = 80'hC089756C6120656C6569;
        inPKT[1162]     = 80'hC08A66656E6420656666;
        inPKT[1163]     = 80'hC08B6963697475722E20;
        inPKT[1164]     = 80'hC08C536564206174206C;
        inPKT[1165]     = 80'hC08D6163757320656C69;
        inPKT[1166]     = 80'hC08E742E205068617365;
        inPKT[1167]     = 80'hC08F6C6C757320656765;
        inPKT[1168]     = 80'hC09074206E6962682076;
        inPKT[1169]     = 80'hC09169746165206D6920;
        inPKT[1170]     = 80'hC0927363656C65726973;
        inPKT[1171]     = 80'hC093717565206665726D;
        inPKT[1172]     = 80'hC094656E74756D207369;
        inPKT[1173]     = 80'hC0957420616D65742076;
        inPKT[1174]     = 80'hC096656C206E65717565;
        inPKT[1175]     = 80'hC0972E204E756E63206C;
        inPKT[1176]     = 80'hC098756374757320616C;
        inPKT[1177]     = 80'hC0996971756574206961;
        inPKT[1178]     = 80'hC09A63756C69732E2050;
        inPKT[1179]     = 80'hC09B72616573656E7420;
        inPKT[1180]     = 80'hC09C6F64696F206A7573;
        inPKT[1181]     = 80'hC09D746F2C20696D7065;
        inPKT[1182]     = 80'hC09E7264696574206E65;
        inPKT[1183]     = 80'hC09F63206C6163757320;
        inPKT[1184]     = 80'hC0A065742C2074656D70;
        inPKT[1185]     = 80'hC0A17573206461706962;
        inPKT[1186]     = 80'hC0A2757320617263752E;
        inPKT[1187]     = 80'hC0A30D0A0D0A43757261;
        inPKT[1188]     = 80'hC0A4626974757220626C;
        inPKT[1189]     = 80'hC0A5616E646974206E75;
        inPKT[1190]     = 80'hC0A66C6C61206964206C;
        inPKT[1191]     = 80'hC0A76F72656D20766F6C;
        inPKT[1192]     = 80'hC0A87574706174206175;
        inPKT[1193]     = 80'hC0A963746F722E204E75;
        inPKT[1194]     = 80'hC0AA6C6C612074696E63;
        inPKT[1195]     = 80'hC0AB6964756E74207465;
        inPKT[1196]     = 80'hC0AC6C6C757320706C61;
        inPKT[1197]     = 80'hC0AD6365726174207075;
        inPKT[1198]     = 80'hC0AE727573206D617869;
        inPKT[1199]     = 80'hC0AF6D757320696D7065;
        inPKT[1200]     = 80'hC0B072646965742E2041;
        inPKT[1201]     = 80'hC0B16C697175616D206E;
        inPKT[1202]     = 80'hC0B26962682074757270;
        inPKT[1203]     = 80'hC0B369732C20616C6971;
        inPKT[1204]     = 80'hC0B475616D2061632076;
        inPKT[1205]     = 80'hC0B5656C69742061632C;
        inPKT[1206]     = 80'hC0B6206D6F6C6C697320;
        inPKT[1207]     = 80'hC0B7736F6C6C69636974;
        inPKT[1208]     = 80'hC0B87564696E206C6962;
        inPKT[1209]     = 80'hC0B965726F2E204D6165;
        inPKT[1210]     = 80'hC0BA63656E6173207075;
        inPKT[1211]     = 80'hC0BB727573206C696775;
        inPKT[1212]     = 80'hC0BC6C612C206C616369;
        inPKT[1213]     = 80'hC0BD6E6961206E656320;
        inPKT[1214]     = 80'hC0BE657820696E2C2075;
        inPKT[1215]     = 80'hC0BF6C6C616D636F7270;
        inPKT[1216]     = 80'hC0C06572207072657469;
        inPKT[1217]     = 80'hC0C1756D20617263752E;
        inPKT[1218]     = 80'hC0C22050656C6C656E74;
        inPKT[1219]     = 80'hC0C36573717565206672;
        inPKT[1220]     = 80'hC0C4696E67696C6C612C;
        inPKT[1221]     = 80'hC0C52065726174207365;
        inPKT[1222]     = 80'hC0C66420666575676961;
        inPKT[1223]     = 80'hC0C77420736167697474;
        inPKT[1224]     = 80'hC0C869732C2061726375;
        inPKT[1225]     = 80'hC0C9206A7573746F2069;
        inPKT[1226]     = 80'hC0CA6E74657264756D20;
        inPKT[1227]     = 80'hC0CB6E6973692C20696E;
        inPKT[1228]     = 80'hC0CC20706F7274746974;
        inPKT[1229]     = 80'hC0CD6F72206D61676E61;
        inPKT[1230]     = 80'hC0CE2076656C69742073;
        inPKT[1231]     = 80'hC0CF65642065782E2053;
        inPKT[1232]     = 80'hC0D0656420617420636F;
        inPKT[1233]     = 80'hC0D16D6D6F646F206572;
        inPKT[1234]     = 80'hC0D26F732C206D6F6C6C;
        inPKT[1235]     = 80'hC0D36973206D61747469;
        inPKT[1236]     = 80'hC0D4732073656D2E204D;
        inPKT[1237]     = 80'hC0D5617572697320656C;
        inPKT[1238]     = 80'hC0D6656D656E74756D20;
        inPKT[1239]     = 80'hC0D76E756E6320736974;
        inPKT[1240]     = 80'hC0D820616D6574206572;
        inPKT[1241]     = 80'hC0D96F7320616363756D;
        inPKT[1242]     = 80'hC0DA73616E2C2076656E;
        inPKT[1243]     = 80'hC0DB656E617469732063;
        inPKT[1244]     = 80'hC0DC6F6E64696D656E74;
        inPKT[1245]     = 80'hC0DD756D206C6967756C;
        inPKT[1246]     = 80'hC0DE612074696E636964;
        inPKT[1247]     = 80'hC0DF756E742E20496E20;
        inPKT[1248]     = 80'hC0E07068617265747261;
        inPKT[1249]     = 80'hC0E120656E696D207268;
        inPKT[1250]     = 80'hC0E26F6E63757320706F;
        inPKT[1251]     = 80'hC0E3737565726520636F;
        inPKT[1252]     = 80'hC0E46E76616C6C69732E;
        inPKT[1253]     = 80'hC0E52043726173206E6F;
        inPKT[1254]     = 80'hC0E66E20657374207665;
        inPKT[1255]     = 80'hC0E76C206C6163757320;
        inPKT[1256]     = 80'hC0E8626C616E64697420;
        inPKT[1257]     = 80'hC0E96D616C6573756164;
        inPKT[1258]     = 80'hC0EA6120637261732061;
        inPKT[1259]     = 80'hC0EB6D65742E00000000;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;
	
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns", countOUT, $time);
	end

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule

