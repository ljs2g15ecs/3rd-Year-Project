`include "SIMON_defintions.svh"

module test_SIMON_3264_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 2400
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 80'hE0001918111009080100;
        inPKT[1]        = 80'hC0014C6F72656D206970;
        inPKT[2]        = 80'hC00273756D20646F6C6F;
        inPKT[3]        = 80'hC003722073697420616D;
        inPKT[4]        = 80'hC00465742C20636F6E73;
        inPKT[5]        = 80'hC0056563746574757220;
        inPKT[6]        = 80'hC0066164697069736369;
        inPKT[7]        = 80'hC0076E6720656C69742E;
        inPKT[8]        = 80'hC0082043757261626974;
        inPKT[9]        = 80'hC009757220756C6C616D;
        inPKT[10]       = 80'hC00A636F727065722074;
        inPKT[11]       = 80'hC00B656D707573206E69;
        inPKT[12]       = 80'hC00C73692C2065742070;
        inPKT[13]       = 80'hC00D6F73756572652075;
        inPKT[14]       = 80'hC00E726E612E2041656E;
        inPKT[15]       = 80'hC00F65616E2073656420;
        inPKT[16]       = 80'hC0106772617669646120;
        inPKT[17]       = 80'hC0116C616375732E204E;
        inPKT[18]       = 80'hC012756C6C6120666163;
        inPKT[19]       = 80'hC013696C6973692E204E;
        inPKT[20]       = 80'hC014756C6C612074656D;
        inPKT[21]       = 80'hC015707573206F726369;
        inPKT[22]       = 80'hC016207175697320656C;
        inPKT[23]       = 80'hC0176974206665756769;
        inPKT[24]       = 80'hC01861742C2076656C20;
        inPKT[25]       = 80'hC01973656D706572206C;
        inPKT[26]       = 80'hC01A656F20696D706572;
        inPKT[27]       = 80'hC01B646965742E204D61;
        inPKT[28]       = 80'hC01C6563656E61732065;
        inPKT[29]       = 80'hC01D74206E756E632069;
        inPKT[30]       = 80'hC01E6E206E6962682066;
        inPKT[31]       = 80'hC01F6163696C69736973;
        inPKT[32]       = 80'hC02020636F6E76616C6C;
        inPKT[33]       = 80'hC02169732E2053656420;
        inPKT[34]       = 80'hC022636F6E6775652068;
        inPKT[35]       = 80'hC023656E647265726974;
        inPKT[36]       = 80'hC02420696163756C6973;
        inPKT[37]       = 80'hC0252E20566976616D75;
        inPKT[38]       = 80'hC0267320766568696375;
        inPKT[39]       = 80'hC0276C61206C75637475;
        inPKT[40]       = 80'hC02873206573742C2076;
        inPKT[41]       = 80'hC0296974616520737573;
        inPKT[42]       = 80'hC02A6369706974206E69;
        inPKT[43]       = 80'hC02B736C20706F727474;
        inPKT[44]       = 80'hC02C69746F722061632E;
        inPKT[45]       = 80'hC02D0D0A0D0A446F6E65;
        inPKT[46]       = 80'hC02E63206D6F6C657374;
        inPKT[47]       = 80'hC02F6965207361706965;
        inPKT[48]       = 80'hC0306E2069642076756C;
        inPKT[49]       = 80'hC0317075746174652076;
        inPKT[50]       = 80'hC0326573746962756C75;
        inPKT[51]       = 80'hC0336D2E204E756C6C61;
        inPKT[52]       = 80'hC03420696E206C696775;
        inPKT[53]       = 80'hC0356C61206672696E67;
        inPKT[54]       = 80'hC036696C6C612C20756C;
        inPKT[55]       = 80'hC0376C616D636F727065;
        inPKT[56]       = 80'hC038722075726E612065;
        inPKT[57]       = 80'hC039742C20706F727474;
        inPKT[58]       = 80'hC03A69746F72206C6563;
        inPKT[59]       = 80'hC03B7475732E20517569;
        inPKT[60]       = 80'hC03C7371756520626C61;
        inPKT[61]       = 80'hC03D6E64697420657520;
        inPKT[62]       = 80'hC03E6D61757269732061;
        inPKT[63]       = 80'hC03F632068656E647265;
        inPKT[64]       = 80'hC0407269742E204E756C;
        inPKT[65]       = 80'hC0416C612076656E656E;
        inPKT[66]       = 80'hC042617469732C206D65;
        inPKT[67]       = 80'hC043747573206574206C;
        inPKT[68]       = 80'hC0447563747573206672;
        inPKT[69]       = 80'hC045696E67696C6C612C;
        inPKT[70]       = 80'hC046206E696268207665;
        inPKT[71]       = 80'hC0476C697420756C6C61;
        inPKT[72]       = 80'hC0486D636F7270657220;
        inPKT[73]       = 80'hC0496469616D2C206567;
        inPKT[74]       = 80'hC04A6574206566666963;
        inPKT[75]       = 80'hC04B6974757220697073;
        inPKT[76]       = 80'hC04C756D207475727069;
        inPKT[77]       = 80'hC04D73206174206E6962;
        inPKT[78]       = 80'hC04E682E205574206567;
        inPKT[79]       = 80'hC04F6574207072657469;
        inPKT[80]       = 80'hC050756D2065726F732C;
        inPKT[81]       = 80'hC0512065676574206469;
        inPKT[82]       = 80'hC0526374756D206C6163;
        inPKT[83]       = 80'hC05375732E204D616563;
        inPKT[84]       = 80'hC054656E617320757420;
        inPKT[85]       = 80'hC055656E696D2065782E;
        inPKT[86]       = 80'hC0562041656E65616E20;
        inPKT[87]       = 80'hC0577669746165207365;
        inPKT[88]       = 80'hC0586D7065722066656C;
        inPKT[89]       = 80'hC05969732C2073656420;
        inPKT[90]       = 80'hC05A756C747269636965;
        inPKT[91]       = 80'hC05B732072697375732E;
        inPKT[92]       = 80'hC05C20446F6E65632063;
        inPKT[93]       = 80'hC05D6F6E736563746574;
        inPKT[94]       = 80'hC05E7572206D69206E69;
        inPKT[95]       = 80'hC05F736C2C2061742063;
        inPKT[96]       = 80'hC0607572737573206970;
        inPKT[97]       = 80'hC06173756D2067726176;
        inPKT[98]       = 80'hC06269646120612E2050;
        inPKT[99]       = 80'hC063686173656C6C7573;
        inPKT[100]      = 80'hC0642073697420616D65;
        inPKT[101]      = 80'hC06574206D61676E6120;
        inPKT[102]      = 80'hC06676656C2069707375;
        inPKT[103]      = 80'hC0676D20656765737461;
        inPKT[104]      = 80'hC0687320706F7274612E;
        inPKT[105]      = 80'hC06920566976616D7573;
        inPKT[106]      = 80'hC06A206C756374757320;
        inPKT[107]      = 80'hC06B656E696D20656765;
        inPKT[108]      = 80'hC06C742074656D706F72;
        inPKT[109]      = 80'hC06D2073616769747469;
        inPKT[110]      = 80'hC06E732E20416C697175;
        inPKT[111]      = 80'hC06F616D20626962656E;
        inPKT[112]      = 80'hC07064756D2073656D20;
        inPKT[113]      = 80'hC0716120636F6E736563;
        inPKT[114]      = 80'hC0727465747572206566;
        inPKT[115]      = 80'hC073666963697475722E;
        inPKT[116]      = 80'hC07420446F6E65632073;
        inPKT[117]      = 80'hC07563656C6572697371;
        inPKT[118]      = 80'hC076756520616C697175;
        inPKT[119]      = 80'hC077616D206375727375;
        inPKT[120]      = 80'hC078732E204375726162;
        inPKT[121]      = 80'hC0796974757220736974;
        inPKT[122]      = 80'hC07A20616D6574206269;
        inPKT[123]      = 80'hC07B62656E64756D2065;
        inPKT[124]      = 80'hC07C6C69742E20536564;
        inPKT[125]      = 80'hC07D206469616D206A75;
        inPKT[126]      = 80'hC07E73746F2C20696163;
        inPKT[127]      = 80'hC07F756C697320717569;
        inPKT[128]      = 80'hC08073206E756C6C6120;
        inPKT[129]      = 80'hC08176697461652C2061;
        inPKT[130]      = 80'hC0826C697175616D2065;
        inPKT[131]      = 80'hC0837569736D6F642066;
        inPKT[132]      = 80'hC084656C69732E0D0A0D;
        inPKT[133]      = 80'hC0850A50726F696E2064;
        inPKT[134]      = 80'hC0866170696275732C20;
        inPKT[135]      = 80'hC0876469616D2076756C;
        inPKT[136]      = 80'hC0887075746174652066;
        inPKT[137]      = 80'hC08972696E67696C6C61;
        inPKT[138]      = 80'hC08A206D616C65737561;
        inPKT[139]      = 80'hC08B64612C206A757374;
        inPKT[140]      = 80'hC08C6F20707572757320;
        inPKT[141]      = 80'hC08D636F6D6D6F646F20;
        inPKT[142]      = 80'hC08E646F6C6F722C2075;
        inPKT[143]      = 80'hC08F742064696374756D;
        inPKT[144]      = 80'hC0902065726174206E75;
        inPKT[145]      = 80'hC0916E63207275747275;
        inPKT[146]      = 80'hC0926D2075726E612E20;
        inPKT[147]      = 80'hC0934E756C6C61206772;
        inPKT[148]      = 80'hC0946176696461207572;
        inPKT[149]      = 80'hC0956E61207669746165;
        inPKT[150]      = 80'hC09620696D7065726469;
        inPKT[151]      = 80'hC0976574206C616F7265;
        inPKT[152]      = 80'hC09865742E2050656C6C;
        inPKT[153]      = 80'hC099656E746573717565;
        inPKT[154]      = 80'hC09A2072686F6E637573;
        inPKT[155]      = 80'hC09B20626962656E6475;
        inPKT[156]      = 80'hC09C6D206E6962682C20;
        inPKT[157]      = 80'hC09D6964206D6F6C6C69;
        inPKT[158]      = 80'hC09E73206469616D2073;
        inPKT[159]      = 80'hC09F7573636970697420;
        inPKT[160]      = 80'hC0A061632E2050656C6C;
        inPKT[161]      = 80'hC0A1656E746573717565;
        inPKT[162]      = 80'hC0A22076656C20696163;
        inPKT[163]      = 80'hC0A3756C697320647569;
        inPKT[164]      = 80'hC0A42E204D6F72626920;
        inPKT[165]      = 80'hC0A5617420616C697175;
        inPKT[166]      = 80'hC0A66574206D61737361;
        inPKT[167]      = 80'hC0A72E2050726F696E20;
        inPKT[168]      = 80'hC0A87669746165206F72;
        inPKT[169]      = 80'hC0A96E617265206F6469;
        inPKT[170]      = 80'hC0AA6F2C206575207675;
        inPKT[171]      = 80'hC0AB6C70757461746520;
        inPKT[172]      = 80'hC0AC697073756D2E2050;
        inPKT[173]      = 80'hC0AD726F696E206C6F62;
        inPKT[174]      = 80'hC0AE6F727469732C2073;
        inPKT[175]      = 80'hC0AF656D206E65632065;
        inPKT[176]      = 80'hC0B07569736D6F642074;
        inPKT[177]      = 80'hC0B1696E636964756E74;
        inPKT[178]      = 80'hC0B22C20617567756520;
        inPKT[179]      = 80'hC0B36D61757269732073;
        inPKT[180]      = 80'hC0B463656C6572697371;
        inPKT[181]      = 80'hC0B57565206D61676E61;
        inPKT[182]      = 80'hC0B62C20657420706F73;
        inPKT[183]      = 80'hC0B775657265206D6920;
        inPKT[184]      = 80'hC0B86E69736C206E6563;
        inPKT[185]      = 80'hC0B9206E6973692E2046;
        inPKT[186]      = 80'hC0BA7573636520656C69;
        inPKT[187]      = 80'hC0BB74206E657175652C;
        inPKT[188]      = 80'hC0BC2076617269757320;
        inPKT[189]      = 80'hC0BD6574206672696E67;
        inPKT[190]      = 80'hC0BE696C6C6120766974;
        inPKT[191]      = 80'hC0BF61652C2076617269;
        inPKT[192]      = 80'hC0C075732076656C206E;
        inPKT[193]      = 80'hC0C1657175652E204E75;
        inPKT[194]      = 80'hC0C26C6C612065742074;
        inPKT[195]      = 80'hC0C3656D707573206A75;
        inPKT[196]      = 80'hC0C473746F2E204D6F72;
        inPKT[197]      = 80'hC0C5626920756C6C616D;
        inPKT[198]      = 80'hC0C6636F727065722073;
        inPKT[199]      = 80'hC0C77573636970697420;
        inPKT[200]      = 80'hC0C8636F6E6775652E20;
        inPKT[201]      = 80'hC0C953656420656C6569;
        inPKT[202]      = 80'hC0CA66656E64206F6469;
        inPKT[203]      = 80'hC0CB6F20616320737573;
        inPKT[204]      = 80'hC0CC6369706974206469;
        inPKT[205]      = 80'hC0CD676E697373696D2E;
        inPKT[206]      = 80'hC0CE2051756973717565;
        inPKT[207]      = 80'hC0CF20616E746520656E;
        inPKT[208]      = 80'hC0D0696D2C20626C616E;
        inPKT[209]      = 80'hC0D164697420696E2063;
        inPKT[210]      = 80'hC0D26F6E736571756174;
        inPKT[211]      = 80'hC0D32061632C20696E74;
        inPKT[212]      = 80'hC0D4657264756D207669;
        inPKT[213]      = 80'hC0D57461652070757275;
        inPKT[214]      = 80'hC0D6732E204D61757269;
        inPKT[215]      = 80'hC0D77320657569736D6F;
        inPKT[216]      = 80'hC0D86420706F73756572;
        inPKT[217]      = 80'hC0D965206C6563747573;
        inPKT[218]      = 80'hC0DA2E20566976616D75;
        inPKT[219]      = 80'hC0DB7320696E74657264;
        inPKT[220]      = 80'hC0DC756D207175616D20;
        inPKT[221]      = 80'hC0DD65752073656D7065;
        inPKT[222]      = 80'hC0DE7220666175636962;
        inPKT[223]      = 80'hC0DF75732E0D0A0D0A49;
        inPKT[224]      = 80'hC0E06E206D6F6C657374;
        inPKT[225]      = 80'hC0E16965206E756C6C61;
        inPKT[226]      = 80'hC0E220616E74652C2061;
        inPKT[227]      = 80'hC0E36320696E74657264;
        inPKT[228]      = 80'hC0E4756D206D61676E61;
        inPKT[229]      = 80'hC0E520636F6E64696D65;
        inPKT[230]      = 80'hC0E66E74756D20636F6E;
        inPKT[231]      = 80'hC0E764696D656E74756D;
        inPKT[232]      = 80'hC0E82E20447569732075;
        inPKT[233]      = 80'hC0E96C74726963696573;
        inPKT[234]      = 80'hC0EA20736F64616C6573;
        inPKT[235]      = 80'hC0EB206E756C6C612C20;
        inPKT[236]      = 80'hC0EC73697420616D6574;
        inPKT[237]      = 80'hC0ED20756C6C616D636F;
        inPKT[238]      = 80'hC0EE72706572206F6469;
        inPKT[239]      = 80'hC0EF6F20707265746975;
        inPKT[240]      = 80'hC0F06D206E65632E2046;
        inPKT[241]      = 80'hC0F17573636520736564;
        inPKT[242]      = 80'hC0F22072697375732070;
        inPKT[243]      = 80'hC0F3656C6C656E746573;
        inPKT[244]      = 80'hC0F47175652C20636F6E;
        inPKT[245]      = 80'hC0F576616C6C69732073;
        inPKT[246]      = 80'hC0F6656D20656765742C;
        inPKT[247]      = 80'hC0F72068656E64726572;
        inPKT[248]      = 80'hC0F8697420657261742E;
        inPKT[249]      = 80'hC0F9204D6F7262692073;
        inPKT[250]      = 80'hC0FA6F64616C65732076;
        inPKT[251]      = 80'hC0FB65686963756C6120;
        inPKT[252]      = 80'hC0FC6C6F626F72746973;
        inPKT[253]      = 80'hC0FD2E2041656E65616E;
        inPKT[254]      = 80'hC0FE206120746F72746F;
        inPKT[255]      = 80'hC0FF7220637572737573;
        inPKT[256]      = 80'hC0002C207363656C6572;
        inPKT[257]      = 80'hC0016973717565206C69;
        inPKT[258]      = 80'hC00267756C6120706F72;
        inPKT[259]      = 80'hC003747469746F722C20;
        inPKT[260]      = 80'hC0046567657374617320;
        inPKT[261]      = 80'hC00565726F732E204475;
        inPKT[262]      = 80'hC00669732074696E6369;
        inPKT[263]      = 80'hC00764756E7420746F72;
        inPKT[264]      = 80'hC008746F722069642070;
        inPKT[265]      = 80'hC0096F73756572652067;
        inPKT[266]      = 80'hC00A7261766964612E20;
        inPKT[267]      = 80'hC00B496E20636F6E7661;
        inPKT[268]      = 80'hC00C6C6C6973206D6920;
        inPKT[269]      = 80'hC00D696420697073756D;
        inPKT[270]      = 80'hC00E206D616C65737561;
        inPKT[271]      = 80'hC00F64612C2075742064;
        inPKT[272]      = 80'hC010696374756D206572;
        inPKT[273]      = 80'hC0116F7320696D706572;
        inPKT[274]      = 80'hC012646965742E205072;
        inPKT[275]      = 80'hC0136F696E20756C6C61;
        inPKT[276]      = 80'hC0146D636F727065722C;
        inPKT[277]      = 80'hC015206D617572697320;
        inPKT[278]      = 80'hC0166964207661726975;
        inPKT[279]      = 80'hC0177320636F6E677565;
        inPKT[280]      = 80'hC0182C2065726F732073;
        inPKT[281]      = 80'hC019617069656E207268;
        inPKT[282]      = 80'hC01A6F6E637573206D69;
        inPKT[283]      = 80'hC01B2C20617420617563;
        inPKT[284]      = 80'hC01C746F72206E657175;
        inPKT[285]      = 80'hC01D652061726375206C;
        inPKT[286]      = 80'hC01E616F726565742064;
        inPKT[287]      = 80'hC01F69616D2E0D0A0D0A;
        inPKT[288]      = 80'hC020467573636520706F;
        inPKT[289]      = 80'hC02172747469746F7220;
        inPKT[290]      = 80'hC0226C696265726F2061;
        inPKT[291]      = 80'hC0237263752C206C6163;
        inPKT[292]      = 80'hC024696E69612068656E;
        inPKT[293]      = 80'hC0256472657269742064;
        inPKT[294]      = 80'hC02669616D20636F6E76;
        inPKT[295]      = 80'hC027616C6C6973207365;
        inPKT[296]      = 80'hC028642E205068617365;
        inPKT[297]      = 80'hC0296C6C7573206E6F6E;
        inPKT[298]      = 80'hC02A2074757270697320;
        inPKT[299]      = 80'hC02B7068617265747261;
        inPKT[300]      = 80'hC02C2C20756C6C616D63;
        inPKT[301]      = 80'hC02D6F72706572206E65;
        inPKT[302]      = 80'hC02E7175652076656C2C;
        inPKT[303]      = 80'hC02F20736F6C6C696369;
        inPKT[304]      = 80'hC030747564696E207665;
        inPKT[305]      = 80'hC0316C69742E2050656C;
        inPKT[306]      = 80'hC0326C656E7465737175;
        inPKT[307]      = 80'hC0336520686162697461;
        inPKT[308]      = 80'hC0346E74206D6F726269;
        inPKT[309]      = 80'hC0352074726973746971;
        inPKT[310]      = 80'hC03675652073656E6563;
        inPKT[311]      = 80'hC037747573206574206E;
        inPKT[312]      = 80'hC0386574757320657420;
        inPKT[313]      = 80'hC0396D616C6573756164;
        inPKT[314]      = 80'hC03A612066616D657320;
        inPKT[315]      = 80'hC03B6163207475727069;
        inPKT[316]      = 80'hC03C7320656765737461;
        inPKT[317]      = 80'hC03D732E204E616D206E;
        inPKT[318]      = 80'hC03E6563207361706965;
        inPKT[319]      = 80'hC03F6E206D6F6C657374;
        inPKT[320]      = 80'hC04069652C2064696374;
        inPKT[321]      = 80'hC041756D206D61737361;
        inPKT[322]      = 80'hC04220656765742C2065;
        inPKT[323]      = 80'hC043676573746173206F;
        inPKT[324]      = 80'hC04464696F2E20457469;
        inPKT[325]      = 80'hC045616D206172637520;
        inPKT[326]      = 80'hC04673617069656E2C20;
        inPKT[327]      = 80'hC0477072657469756D20;
        inPKT[328]      = 80'hC04861206D6F6C6C6973;
        inPKT[329]      = 80'hC04920612C2076756C70;
        inPKT[330]      = 80'hC04A7574617465206E6F;
        inPKT[331]      = 80'hC04B6E20657261742E20;
        inPKT[332]      = 80'hC04C5574207669746165;
        inPKT[333]      = 80'hC04D206E696268206C6F;
        inPKT[334]      = 80'hC04E626F72746973206C;
        inPKT[335]      = 80'hC04F6563747573206661;
        inPKT[336]      = 80'hC0507563696275732070;
        inPKT[337]      = 80'hC0516F72746120657520;
        inPKT[338]      = 80'hC05273697420616D6574;
        inPKT[339]      = 80'hC053206E69736C2E204D;
        inPKT[340]      = 80'hC0546F72626920706F72;
        inPKT[341]      = 80'hC055747469746F722076;
        inPKT[342]      = 80'hC056656C697420657520;
        inPKT[343]      = 80'hC057646F6C6F72206C61;
        inPKT[344]      = 80'hC0586F726565742C2073;
        inPKT[345]      = 80'hC059697420616D657420;
        inPKT[346]      = 80'hC05A696D706572646965;
        inPKT[347]      = 80'hC05B7420656E696D2073;
        inPKT[348]      = 80'hC05C6F64616C65732E20;
        inPKT[349]      = 80'hC05D4E756C6C616D2075;
        inPKT[350]      = 80'hC05E6C6C616D636F7270;
        inPKT[351]      = 80'hC05F6572207475727069;
        inPKT[352]      = 80'hC060732061742070656C;
        inPKT[353]      = 80'hC0616C656E7465737175;
        inPKT[354]      = 80'hC0626520766172697573;
        inPKT[355]      = 80'hC0632E20566976616D75;
        inPKT[356]      = 80'hC0647320657520696D70;
        inPKT[357]      = 80'hC065657264696574206E;
        inPKT[358]      = 80'hC066657175652E205365;
        inPKT[359]      = 80'hC0676420717569732061;
        inPKT[360]      = 80'hC0687563746F7220616E;
        inPKT[361]      = 80'hC06974652E204D617572;
        inPKT[362]      = 80'hC06A69732073656D7065;
        inPKT[363]      = 80'hC06B7220697073756D20;
        inPKT[364]      = 80'hC06C7365642064756920;
        inPKT[365]      = 80'hC06D706F73756572652C;
        inPKT[366]      = 80'hC06E20617420616C6971;
        inPKT[367]      = 80'hC06F75616D206D657475;
        inPKT[368]      = 80'hC0707320656C65696665;
        inPKT[369]      = 80'hC0716E642E204E756C6C;
        inPKT[370]      = 80'hC072616D207472697374;
        inPKT[371]      = 80'hC0736971756520656C65;
        inPKT[372]      = 80'hC0746966656E64206572;
        inPKT[373]      = 80'hC0756F732C2065676574;
        inPKT[374]      = 80'hC076206665726D656E74;
        inPKT[375]      = 80'hC077756D20697073756D;
        inPKT[376]      = 80'hC07820656C656D656E74;
        inPKT[377]      = 80'hC079756D206E65632E0D;
        inPKT[378]      = 80'hC07A0A0D0A50656C6C65;
        inPKT[379]      = 80'hC07B6E74657371756520;
        inPKT[380]      = 80'hC07C68656E6472657269;
        inPKT[381]      = 80'hC07D7420626962656E64;
        inPKT[382]      = 80'hC07E756D206C6967756C;
        inPKT[383]      = 80'hC07F612C20657420736F;
        inPKT[384]      = 80'hC08064616C6573206D61;
        inPKT[385]      = 80'hC081676E612064617069;
        inPKT[386]      = 80'hC08262757320696E2E20;
        inPKT[387]      = 80'hC083496E20616C697175;
        inPKT[388]      = 80'hC084657420746F72746F;
        inPKT[389]      = 80'hC0857220656765742063;
        inPKT[390]      = 80'hC0866F6E736563746574;
        inPKT[391]      = 80'hC087757220636F6E7365;
        inPKT[392]      = 80'hC0886374657475722E20;
        inPKT[393]      = 80'hC0895175697371756520;
        inPKT[394]      = 80'hC08A7472697374697175;
        inPKT[395]      = 80'hC08B6520726973757320;
        inPKT[396]      = 80'hC08C657261742C206574;
        inPKT[397]      = 80'hC08D20616C6971756574;
        inPKT[398]      = 80'hC08E20656C697420616C;
        inPKT[399]      = 80'hC08F6971756574206575;
        inPKT[400]      = 80'hC0902E20496E74656765;
        inPKT[401]      = 80'hC09172206E6F6E206D61;
        inPKT[402]      = 80'hC092676E6120696E2066;
        inPKT[403]      = 80'hC093656C697320706F72;
        inPKT[404]      = 80'hC094747469746F722073;
        inPKT[405]      = 80'hC095616769747469732E;
        inPKT[406]      = 80'hC0962051756973717565;
        inPKT[407]      = 80'hC0972076697665727261;
        inPKT[408]      = 80'hC098206F726369206163;
        inPKT[409]      = 80'hC0992072757472756D20;
        inPKT[410]      = 80'hC09A6C616F726565742E;
        inPKT[411]      = 80'hC09B2041656E65616E20;
        inPKT[412]      = 80'hC09C636F6E76616C6C69;
        inPKT[413]      = 80'hC09D732064696374756D;
        inPKT[414]      = 80'hC09E207475727069732C;
        inPKT[415]      = 80'hC09F2065742066696E69;
        inPKT[416]      = 80'hC0A06275732073617069;
        inPKT[417]      = 80'hC0A1656E20636F6E6775;
        inPKT[418]      = 80'hC0A26520696E2E205365;
        inPKT[419]      = 80'hC0A36420612065726174;
        inPKT[420]      = 80'hC0A4206F726E6172652C;
        inPKT[421]      = 80'hC0A5206D6F6C6C697320;
        inPKT[422]      = 80'hC0A66E69736C2061632C;
        inPKT[423]      = 80'hC0A7206469676E697373;
        inPKT[424]      = 80'hC0A8696D206E65717565;
        inPKT[425]      = 80'hC0A92E20517569737175;
        inPKT[426]      = 80'hC0AA65206D616C657375;
        inPKT[427]      = 80'hC0AB61646120706F7375;
        inPKT[428]      = 80'hC0AC6572652074757270;
        inPKT[429]      = 80'hC0AD697320657520756C;
        inPKT[430]      = 80'hC0AE6C616D636F727065;
        inPKT[431]      = 80'hC0AF722E20446F6E6563;
        inPKT[432]      = 80'hC0B02076697665727261;
        inPKT[433]      = 80'hC0B120626962656E6475;
        inPKT[434]      = 80'hC0B26D206E756E632C20;
        inPKT[435]      = 80'hC0B364696374756D2069;
        inPKT[436]      = 80'hC0B46D70657264696574;
        inPKT[437]      = 80'hC0B5206E65717565206D;
        inPKT[438]      = 80'hC0B66178696D75732069;
        inPKT[439]      = 80'hC0B76E2E20446F6E6563;
        inPKT[440]      = 80'hC0B820757420756C7472;
        inPKT[441]      = 80'hC0B96963657320646F6C;
        inPKT[442]      = 80'hC0BA6F722E2056697661;
        inPKT[443]      = 80'hC0BB6D75732073656420;
        inPKT[444]      = 80'hC0BC6175677565207072;
        inPKT[445]      = 80'hC0BD657469756D2C2076;
        inPKT[446]      = 80'hC0BE6F6C757470617420;
        inPKT[447]      = 80'hC0BF657261742061632C;
        inPKT[448]      = 80'hC0C020706F7274612064;
        inPKT[449]      = 80'hC0C169616D2E204D6175;
        inPKT[450]      = 80'hC0C272697320696E2070;
        inPKT[451]      = 80'hC0C37572757320756C74;
        inPKT[452]      = 80'hC0C47269636965732C20;
        inPKT[453]      = 80'hC0C57375736369706974;
        inPKT[454]      = 80'hC0C6206469616D207365;
        inPKT[455]      = 80'hC0C7642C2074696E6369;
        inPKT[456]      = 80'hC0C864756E7420656E69;
        inPKT[457]      = 80'hC0C96D2E20446F6E6563;
        inPKT[458]      = 80'hC0CA207175697320706F;
        inPKT[459]      = 80'hC0CB7375657265206E69;
        inPKT[460]      = 80'hC0CC62682E20496E2068;
        inPKT[461]      = 80'hC0CD6163206861626974;
        inPKT[462]      = 80'hC0CE6173736520706C61;
        inPKT[463]      = 80'hC0CF7465612064696374;
        inPKT[464]      = 80'hC0D0756D73742E0D0A0D;
        inPKT[465]      = 80'hC0D10A4D6F726269206F;
        inPKT[466]      = 80'hC0D2726E617265206A75;
        inPKT[467]      = 80'hC0D373746F2061742071;
        inPKT[468]      = 80'hC0D475616D2066617563;
        inPKT[469]      = 80'hC0D5696275732C207369;
        inPKT[470]      = 80'hC0D67420616D6574206D;
        inPKT[471]      = 80'hC0D76F6C657374696520;
        inPKT[472]      = 80'hC0D86C656F2063757273;
        inPKT[473]      = 80'hC0D975732E204D617572;
        inPKT[474]      = 80'hC0DA6973206C616F7265;
        inPKT[475]      = 80'hC0DB657420616E746520;
        inPKT[476]      = 80'hC0DC61206D6574757320;
        inPKT[477]      = 80'hC0DD6566666963697475;
        inPKT[478]      = 80'hC0DE7220766172697573;
        inPKT[479]      = 80'hC0DF2E20536564207665;
        inPKT[480]      = 80'hC0E06C206F7263692073;
        inPKT[481]      = 80'hC0E16167697474697320;
        inPKT[482]      = 80'hC0E26E756E6320626C61;
        inPKT[483]      = 80'hC0E36E64697420636F6E;
        inPKT[484]      = 80'hC0E47365717561742E20;
        inPKT[485]      = 80'hC0E55072616573656E74;
        inPKT[486]      = 80'hC0E6206D616C65737561;
        inPKT[487]      = 80'hC0E76461206E65717565;
        inPKT[488]      = 80'hC0E82071756973206469;
        inPKT[489]      = 80'hC0E96374756D20646967;
        inPKT[490]      = 80'hC0EA6E697373696D2E20;
        inPKT[491]      = 80'hC0EB446F6E6563206661;
        inPKT[492]      = 80'hC0EC63696C6973697320;
        inPKT[493]      = 80'hC0ED73697420616D6574;
        inPKT[494]      = 80'hC0EE2076656C69742065;
        inPKT[495]      = 80'hC0EF75206C6F626F7274;
        inPKT[496]      = 80'hC0F069732E204E756C6C;
        inPKT[497]      = 80'hC0F1616D20626C616E64;
        inPKT[498]      = 80'hC0F2697420656C656D65;
        inPKT[499]      = 80'hC0F36E74756D206D6175;
        inPKT[500]      = 80'hC0F47269732C20766974;
        inPKT[501]      = 80'hC0F5616520656C656D65;
        inPKT[502]      = 80'hC0F66E74756D20646F6C;
        inPKT[503]      = 80'hC0F76F722068656E6472;
        inPKT[504]      = 80'hC0F86572697420766974;
        inPKT[505]      = 80'hC0F961652E2046757363;
        inPKT[506]      = 80'hC0FA65206D6F6C657374;
        inPKT[507]      = 80'hC0FB69652C20656C6974;
        inPKT[508]      = 80'hC0FC20757420616C6971;
        inPKT[509]      = 80'hC0FD75657420766F6C75;
        inPKT[510]      = 80'hC0FE747061742C206E65;
        inPKT[511]      = 80'hC0FF7175652076656C69;
        inPKT[512]      = 80'hC0007420707265746975;
        inPKT[513]      = 80'hC0016D2061756775652C;
        inPKT[514]      = 80'hC002206672696E67696C;
        inPKT[515]      = 80'hC0036C6120636F6E6469;
        inPKT[516]      = 80'hC0046D656E74756D206A;
        inPKT[517]      = 80'hC0057573746F20736170;
        inPKT[518]      = 80'hC00669656E2061206A75;
        inPKT[519]      = 80'hC00773746F2E20506861;
        inPKT[520]      = 80'hC00873656C6C75732071;
        inPKT[521]      = 80'hC0097569732061756374;
        inPKT[522]      = 80'hC00A6F72206C6F72656D;
        inPKT[523]      = 80'hC00B2C20696E20616C69;
        inPKT[524]      = 80'hC00C7175616D206E756E;
        inPKT[525]      = 80'hC00D632E20557420656C;
        inPKT[526]      = 80'hC00E656966656E642061;
        inPKT[527]      = 80'hC00F6E7465206574206E;
        inPKT[528]      = 80'hC010697369206D6F6C65;
        inPKT[529]      = 80'hC0117374696520636F6E;
        inPKT[530]      = 80'hC01276616C6C69732069;
        inPKT[531]      = 80'hC013642065742073656D;
        inPKT[532]      = 80'hC0142E20536564206163;
        inPKT[533]      = 80'hC01520626962656E6475;
        inPKT[534]      = 80'hC0166D20617263752E20;
        inPKT[535]      = 80'hC0174675736365207665;
        inPKT[536]      = 80'hC01873746962756C756D;
        inPKT[537]      = 80'hC019206E756E63206567;
        inPKT[538]      = 80'hC01A65742074656C6C75;
        inPKT[539]      = 80'hC01B73206665726D656E;
        inPKT[540]      = 80'hC01C74756D2C206E6563;
        inPKT[541]      = 80'hC01D2072686F6E637573;
        inPKT[542]      = 80'hC01E206D617373612063;
        inPKT[543]      = 80'hC01F6F6D6D6F646F2E20;
        inPKT[544]      = 80'hC0204D616563656E6173;
        inPKT[545]      = 80'hC021206964206E756E63;
        inPKT[546]      = 80'hC022206E6F6E20657820;
        inPKT[547]      = 80'hC023766573746962756C;
        inPKT[548]      = 80'hC024756D206F726E6172;
        inPKT[549]      = 80'hC02565207574206E6563;
        inPKT[550]      = 80'hC0262065726F732E2041;
        inPKT[551]      = 80'hC0276C697175616D2065;
        inPKT[552]      = 80'hC0286666696369747572;
        inPKT[553]      = 80'hC02920636F6D6D6F646F;
        inPKT[554]      = 80'hC02A206469616D206964;
        inPKT[555]      = 80'hC02B206C6F626F727469;
        inPKT[556]      = 80'hC02C732E205365642061;
        inPKT[557]      = 80'hC02D632074656D706F72;
        inPKT[558]      = 80'hC02E206C65637475732E;
        inPKT[559]      = 80'hC02F204E756E6320656C;
        inPKT[560]      = 80'hC030656D656E74756D20;
        inPKT[561]      = 80'hC0317574206C65637475;
        inPKT[562]      = 80'hC032732061632074696E;
        inPKT[563]      = 80'hC033636964756E742E20;
        inPKT[564]      = 80'hC034557420696163756C;
        inPKT[565]      = 80'hC0356973206E756C6C61;
        inPKT[566]      = 80'hC0362071756973206578;
        inPKT[567]      = 80'hC03720656C656D656E74;
        inPKT[568]      = 80'hC038756D2C20616C6971;
        inPKT[569]      = 80'hC0397565742073656D70;
        inPKT[570]      = 80'hC03A6572206D61676E61;
        inPKT[571]      = 80'hC03B20656C656966656E;
        inPKT[572]      = 80'hC03C642E0D0A0D0A4375;
        inPKT[573]      = 80'hC03D7261626974757220;
        inPKT[574]      = 80'hC03E746F72746F72206E;
        inPKT[575]      = 80'hC03F69736C2C20756C74;
        inPKT[576]      = 80'hC0407269636965732069;
        inPKT[577]      = 80'hC0416E206E6571756520;
        inPKT[578]      = 80'hC04261632C2061636375;
        inPKT[579]      = 80'hC0436D73616E20636F6E;
        inPKT[580]      = 80'hC044736571756174206D;
        inPKT[581]      = 80'hC045657475732E204D61;
        inPKT[582]      = 80'hC0466563656E6173206D;
        inPKT[583]      = 80'hC0476173736120736170;
        inPKT[584]      = 80'hC04869656E2C206D6174;
        inPKT[585]      = 80'hC04974697320696E2076;
        inPKT[586]      = 80'hC04A656E656E61746973;
        inPKT[587]      = 80'hC04B2073697420616D65;
        inPKT[588]      = 80'hC04C742C20617563746F;
        inPKT[589]      = 80'hC04D722073697420616D;
        inPKT[590]      = 80'hC04E657420656E696D2E;
        inPKT[591]      = 80'hC04F204E756E63207669;
        inPKT[592]      = 80'hC050746165206D657475;
        inPKT[593]      = 80'hC0517320636F6D6D6F64;
        inPKT[594]      = 80'hC0526F2C206D61747469;
        inPKT[595]      = 80'hC05373206D6173736120;
        inPKT[596]      = 80'hC05473697420616D6574;
        inPKT[597]      = 80'hC0552C20766172697573;
        inPKT[598]      = 80'hC056206C6F72656D2E20;
        inPKT[599]      = 80'hC0574E756E6320696E20;
        inPKT[600]      = 80'hC058656C697420656C69;
        inPKT[601]      = 80'hC059742E204E756E6320;
        inPKT[602]      = 80'hC05A6F726E6172652063;
        inPKT[603]      = 80'hC05B6F6E736563746574;
        inPKT[604]      = 80'hC05C7572206D61676E61;
        inPKT[605]      = 80'hC05D2C2073697420616D;
        inPKT[606]      = 80'hC05E657420706F727474;
        inPKT[607]      = 80'hC05F69746F7220617263;
        inPKT[608]      = 80'hC060752072686F6E6375;
        inPKT[609]      = 80'hC061732065752E205375;
        inPKT[610]      = 80'hC0627370656E64697373;
        inPKT[611]      = 80'hC06365207363656C6572;
        inPKT[612]      = 80'hC064697371756520756C;
        inPKT[613]      = 80'hC0657472696369657320;
        inPKT[614]      = 80'hC0666578206120616C69;
        inPKT[615]      = 80'hC0677175616D2E205375;
        inPKT[616]      = 80'hC0687370656E64697373;
        inPKT[617]      = 80'hC069652072757472756D;
        inPKT[618]      = 80'hC06A20736F6C6C696369;
        inPKT[619]      = 80'hC06B747564696E206E75;
        inPKT[620]      = 80'hC06C6E632C206E6F6E20;
        inPKT[621]      = 80'hC06D636F6E76616C6C69;
        inPKT[622]      = 80'hC06E7320747572706973;
        inPKT[623]      = 80'hC06F206C616F72656574;
        inPKT[624]      = 80'hC0702073697420616D65;
        inPKT[625]      = 80'hC071742E2041656E6561;
        inPKT[626]      = 80'hC0726E20612066696E69;
        inPKT[627]      = 80'hC073627573206D617572;
        inPKT[628]      = 80'hC07469732C2071756973;
        inPKT[629]      = 80'hC0752063757273757320;
        inPKT[630]      = 80'hC0766E756E632E20496E;
        inPKT[631]      = 80'hC0772066657567696174;
        inPKT[632]      = 80'hC078206475692076656C;
        inPKT[633]      = 80'hC0792075726E61207365;
        inPKT[634]      = 80'hC07A6D70657220666175;
        inPKT[635]      = 80'hC07B63696275732E204D;
        inPKT[636]      = 80'hC07C617572697320756C;
        inPKT[637]      = 80'hC07D7472696369657320;
        inPKT[638]      = 80'hC07E6174207475727069;
        inPKT[639]      = 80'hC07F7320656765742070;
        inPKT[640]      = 80'hC080656C6C656E746573;
        inPKT[641]      = 80'hC0817175652E20507261;
        inPKT[642]      = 80'hC0826573656E74207369;
        inPKT[643]      = 80'hC0837420616D6574206C;
        inPKT[644]      = 80'hC0846967756C6120636F;
        inPKT[645]      = 80'hC0856E76616C6C69732C;
        inPKT[646]      = 80'hC08620656C656D656E74;
        inPKT[647]      = 80'hC087756D206E756C6C61;
        inPKT[648]      = 80'hC08820756C6C616D636F;
        inPKT[649]      = 80'hC089727065722C20616C;
        inPKT[650]      = 80'hC08A697175616D207572;
        inPKT[651]      = 80'hC08B6E612E2045746961;
        inPKT[652]      = 80'hC08C6D207175616D2065;
        inPKT[653]      = 80'hC08D6C69742C20706F73;
        inPKT[654]      = 80'hC08E7565726520757420;
        inPKT[655]      = 80'hC08F7175616D20656765;
        inPKT[656]      = 80'hC090742C2066696E6962;
        inPKT[657]      = 80'hC091757320736F6C6C69;
        inPKT[658]      = 80'hC0926369747564696E20;
        inPKT[659]      = 80'hC0936E756C6C612E2049;
        inPKT[660]      = 80'hC0946E20737573636970;
        inPKT[661]      = 80'hC095697420656E696D20;
        inPKT[662]      = 80'hC09665742065726F7320;
        inPKT[663]      = 80'hC09766696E696275732C;
        inPKT[664]      = 80'hC098207574207363656C;
        inPKT[665]      = 80'hC0996572697371756520;
        inPKT[666]      = 80'hC09A74656C6C75732066;
        inPKT[667]      = 80'hC09B6575676961742E20;
        inPKT[668]      = 80'hC09C4375726162697475;
        inPKT[669]      = 80'hC09D72206E6F6E206D61;
        inPKT[670]      = 80'hC09E7373612076617269;
        inPKT[671]      = 80'hC09F757320646F6C6F72;
        inPKT[672]      = 80'hC0A02067726176696461;
        inPKT[673]      = 80'hC0A120656C656D656E74;
        inPKT[674]      = 80'hC0A2756D207175697320;
        inPKT[675]      = 80'hC0A375742066656C6973;
        inPKT[676]      = 80'hC0A42E2050686173656C;
        inPKT[677]      = 80'hC0A56C75732065756973;
        inPKT[678]      = 80'hC0A66D6F642069707375;
        inPKT[679]      = 80'hC0A76D20656765742076;
        inPKT[680]      = 80'hC0A8656C6974206C6F62;
        inPKT[681]      = 80'hC0A96F727469732C2065;
        inPKT[682]      = 80'hC0AA67657420706F7274;
        inPKT[683]      = 80'hC0AB61206D6175726973;
        inPKT[684]      = 80'hC0AC2074656D7075732E;
        inPKT[685]      = 80'hC0AD2053656420696D70;
        inPKT[686]      = 80'hC0AE6572646965742076;
        inPKT[687]      = 80'hC0AF6F6C757470617420;
        inPKT[688]      = 80'hC0B074656C6C75732065;
        inPKT[689]      = 80'hC0B1752074696E636964;
        inPKT[690]      = 80'hC0B2756E742E0D0A0D0A;
        inPKT[691]      = 80'hC0B355742076656C206D;
        inPKT[692]      = 80'hC0B469206174206D6574;
        inPKT[693]      = 80'hC0B57573206672696E67;
        inPKT[694]      = 80'hC0B6696C6C6120677261;
        inPKT[695]      = 80'hC0B7766964612E205072;
        inPKT[696]      = 80'hC0B8616573656E742065;
        inPKT[697]      = 80'hC0B9726F73206E696268;
        inPKT[698]      = 80'hC0BA2C20637572737573;
        inPKT[699]      = 80'hC0BB2065676573746173;
        inPKT[700]      = 80'hC0BC2074696E63696475;
        inPKT[701]      = 80'hC0BD6E7420736F64616C;
        inPKT[702]      = 80'hC0BE65732C207363656C;
        inPKT[703]      = 80'hC0BF6572697371756520;
        inPKT[704]      = 80'hC0C06E65632066656C69;
        inPKT[705]      = 80'hC0C1732E20496E746567;
        inPKT[706]      = 80'hC0C2657220696D706572;
        inPKT[707]      = 80'hC0C364696574206D616C;
        inPKT[708]      = 80'hC0C4657375616461206E;
        inPKT[709]      = 80'hC0C569736C20616C6971;
        inPKT[710]      = 80'hC0C67565742076656E65;
        inPKT[711]      = 80'hC0C76E617469732E2049;
        inPKT[712]      = 80'hC0C86E74656765722073;
        inPKT[713]      = 80'hC0C9656420706F727474;
        inPKT[714]      = 80'hC0CA69746F7220697073;
        inPKT[715]      = 80'hC0CB756D2E20496E7465;
        inPKT[716]      = 80'hC0CC67657220636F6D6D;
        inPKT[717]      = 80'hC0CD6F646F2066657567;
        inPKT[718]      = 80'hC0CE69617420746F7274;
        inPKT[719]      = 80'hC0CF6F722C206575206C;
        inPKT[720]      = 80'hC0D06F626F7274697320;
        inPKT[721]      = 80'hC0D1617567756520656C;
        inPKT[722]      = 80'hC0D2656D656E74756D20;
        inPKT[723]      = 80'hC0D373697420616D6574;
        inPKT[724]      = 80'hC0D42E20446F6E656320;
        inPKT[725]      = 80'hC0D5766573746962756C;
        inPKT[726]      = 80'hC0D6756D206C6967756C;
        inPKT[727]      = 80'hC0D7612061756775652C;
        inPKT[728]      = 80'hC0D82065742066696E69;
        inPKT[729]      = 80'hC0D96275732061726375;
        inPKT[730]      = 80'hC0DA20706F7274612069;
        inPKT[731]      = 80'hC0DB6E2E204E756C6C61;
        inPKT[732]      = 80'hC0DC2073656D2074656C;
        inPKT[733]      = 80'hC0DD6C75732C20756C6C;
        inPKT[734]      = 80'hC0DE616D636F72706572;
        inPKT[735]      = 80'hC0DF2061742063757273;
        inPKT[736]      = 80'hC0E0757320612C20706F;
        inPKT[737]      = 80'hC0E17274612073697420;
        inPKT[738]      = 80'hC0E2616D6574206D6167;
        inPKT[739]      = 80'hC0E36E612E204E756E63;
        inPKT[740]      = 80'hC0E42076697461652069;
        inPKT[741]      = 80'hC0E56D70657264696574;
        inPKT[742]      = 80'hC0E62070757275732C20;
        inPKT[743]      = 80'hC0E76E656320736F6C6C;
        inPKT[744]      = 80'hC0E8696369747564696E;
        inPKT[745]      = 80'hC0E92074656C6C75732E;
        inPKT[746]      = 80'hC0EA20416C697175616D;
        inPKT[747]      = 80'hC0EB206572617420766F;
        inPKT[748]      = 80'hC0EC6C75747061742E20;
        inPKT[749]      = 80'hC0ED536564206964206D;
        inPKT[750]      = 80'hC0EE61676E6120636F6D;
        inPKT[751]      = 80'hC0EF6D6F646F2C206C75;
        inPKT[752]      = 80'hC0F0637475732076656C;
        inPKT[753]      = 80'hC0F1697420717569732C;
        inPKT[754]      = 80'hC0F220657569736D6F64;
        inPKT[755]      = 80'hC0F320656E696D2E2049;
        inPKT[756]      = 80'hC0F46E7465676572206D;
        inPKT[757]      = 80'hC0F5617474697320736F;
        inPKT[758]      = 80'hC0F664616C6573206665;
        inPKT[759]      = 80'hC0F7726D656E74756D2E;
        inPKT[760]      = 80'hC0F82051756973717565;
        inPKT[761]      = 80'hC0F92073656420667269;
        inPKT[762]      = 80'hC0FA6E67696C6C61206C;
        inPKT[763]      = 80'hC0FB6F72656D2E204372;
        inPKT[764]      = 80'hC0FC6173207665686963;
        inPKT[765]      = 80'hC0FD756C612074656D70;
        inPKT[766]      = 80'hC0FE7573207361706965;
        inPKT[767]      = 80'hC0FF6E20757420636F6E;
        inPKT[768]      = 80'hC0006775652E20447569;
        inPKT[769]      = 80'hC001732073617069656E;
        inPKT[770]      = 80'hC00220656E696D2C2070;
        inPKT[771]      = 80'hC0036F727461206E6563;
        inPKT[772]      = 80'hC004206C656F2069642C;
        inPKT[773]      = 80'hC0052065666669636974;
        inPKT[774]      = 80'hC006757220706F737565;
        inPKT[775]      = 80'hC0077265206C69626572;
        inPKT[776]      = 80'hC0086F2E204E756C6C61;
        inPKT[777]      = 80'hC0096D2061632074656D;
        inPKT[778]      = 80'hC00A706F72206D657475;
        inPKT[779]      = 80'hC00B732E205365642076;
        inPKT[780]      = 80'hC00C656C207475727069;
        inPKT[781]      = 80'hC00D7320666575676961;
        inPKT[782]      = 80'hC00E742C20696163756C;
        inPKT[783]      = 80'hC00F6973206175677565;
        inPKT[784]      = 80'hC01020717569732C2074;
        inPKT[785]      = 80'hC011696E636964756E74;
        inPKT[786]      = 80'hC012207475727069732E;
        inPKT[787]      = 80'hC0130D0A0D0A56697661;
        inPKT[788]      = 80'hC0146D757320706F7375;
        inPKT[789]      = 80'hC01565726520706F7274;
        inPKT[790]      = 80'hC0167469746F72206175;
        inPKT[791]      = 80'hC0176775652C20766172;
        inPKT[792]      = 80'hC0186975732061636375;
        inPKT[793]      = 80'hC0196D73616E20656C69;
        inPKT[794]      = 80'hC01A742076756C707574;
        inPKT[795]      = 80'hC01B6174652065676574;
        inPKT[796]      = 80'hC01C2E20517569737175;
        inPKT[797]      = 80'hC01D6520736564206D61;
        inPKT[798]      = 80'hC01E6C65737561646120;
        inPKT[799]      = 80'hC01F6E69736C2E20496E;
        inPKT[800]      = 80'hC02074657264756D2065;
        inPKT[801]      = 80'hC02174206D616C657375;
        inPKT[802]      = 80'hC0226164612066616D65;
        inPKT[803]      = 80'hC0237320616320616E74;
        inPKT[804]      = 80'hC0246520697073756D20;
        inPKT[805]      = 80'hC0257072696D69732069;
        inPKT[806]      = 80'hC0266E20666175636962;
        inPKT[807]      = 80'hC02775732E204E756E63;
        inPKT[808]      = 80'hC0282074757270697320;
        inPKT[809]      = 80'hC0296469616D2C207375;
        inPKT[810]      = 80'hC02A7363697069742061;
        inPKT[811]      = 80'hC02B632065726F732076;
        inPKT[812]      = 80'hC02C656C2C2074656D70;
        inPKT[813]      = 80'hC02D75732076656E656E;
        inPKT[814]      = 80'hC02E6174697320697073;
        inPKT[815]      = 80'hC02F756D2E2044756973;
        inPKT[816]      = 80'hC030206C756374757320;
        inPKT[817]      = 80'hC03172686F6E63757320;
        inPKT[818]      = 80'hC0326D617373612E2046;
        inPKT[819]      = 80'hC0337573636520757420;
        inPKT[820]      = 80'hC0346C6163696E696120;
        inPKT[821]      = 80'hC0357475727069732E20;
        inPKT[822]      = 80'hC036566976616D757320;
        inPKT[823]      = 80'hC03772757472756D2074;
        inPKT[824]      = 80'hC038656C6C7573206175;
        inPKT[825]      = 80'hC0396775652C20617420;
        inPKT[826]      = 80'hC03A6F726E617265206E;
        inPKT[827]      = 80'hC03B69736C2066616369;
        inPKT[828]      = 80'hC03C6C69736973206574;
        inPKT[829]      = 80'hC03D2E204E756E632073;
        inPKT[830]      = 80'hC03E6564206E69736920;
        inPKT[831]      = 80'hC03F72697375732E2049;
        inPKT[832]      = 80'hC0406E74656765722065;
        inPKT[833]      = 80'hC0416C656D656E74756D;
        inPKT[834]      = 80'hC042206D617572697320;
        inPKT[835]      = 80'hC0437175616D2C207574;
        inPKT[836]      = 80'hC044207665686963756C;
        inPKT[837]      = 80'hC04561206D6175726973;
        inPKT[838]      = 80'hC04620636F6E67756520;
        inPKT[839]      = 80'hC04765752E0D0A0D0A46;
        inPKT[840]      = 80'hC0487573636520612074;
        inPKT[841]      = 80'hC049656C6C7573207369;
        inPKT[842]      = 80'hC04A7420616D65742065;
        inPKT[843]      = 80'hC04B726174206665726D;
        inPKT[844]      = 80'hC04C656E74756D207363;
        inPKT[845]      = 80'hC04D656C657269737175;
        inPKT[846]      = 80'hC04E652E204375726162;
        inPKT[847]      = 80'hC04F6974757220696E20;
        inPKT[848]      = 80'hC05076656C6974206174;
        inPKT[849]      = 80'hC05120656E696D206C61;
        inPKT[850]      = 80'hC05263696E6961207665;
        inPKT[851]      = 80'hC053686963756C612061;
        inPKT[852]      = 80'hC05463206964206A7573;
        inPKT[853]      = 80'hC055746F2E2050726F69;
        inPKT[854]      = 80'hC0566E206E6F6E20646F;
        inPKT[855]      = 80'hC0576C6F722065666669;
        inPKT[856]      = 80'hC05863697475722C2074;
        inPKT[857]      = 80'hC059696E636964756E74;
        inPKT[858]      = 80'hC05A206F64696F206575;
        inPKT[859]      = 80'hC05B2C20666175636962;
        inPKT[860]      = 80'hC05C757320656E696D2E;
        inPKT[861]      = 80'hC05D2050656C6C656E74;
        inPKT[862]      = 80'hC05E6573717565206461;
        inPKT[863]      = 80'hC05F7069627573206F72;
        inPKT[864]      = 80'hC0606369206163206C6F;
        inPKT[865]      = 80'hC06172656D2069616375;
        inPKT[866]      = 80'hC0626C69732C20736974;
        inPKT[867]      = 80'hC06320616D657420626C;
        inPKT[868]      = 80'hC064616E646974206172;
        inPKT[869]      = 80'hC0656375207472697374;
        inPKT[870]      = 80'hC066697175652E204165;
        inPKT[871]      = 80'hC0676E65616E20747269;
        inPKT[872]      = 80'hC0687374697175652074;
        inPKT[873]      = 80'hC0696F72746F72206E65;
        inPKT[874]      = 80'hC06A63206A7573746F20;
        inPKT[875]      = 80'hC06B616C697175616D2C;
        inPKT[876]      = 80'hC06C20696E2070726574;
        inPKT[877]      = 80'hC06D69756D2066656C69;
        inPKT[878]      = 80'hC06E73206D6F6C657374;
        inPKT[879]      = 80'hC06F69652E2053656420;
        inPKT[880]      = 80'hC07065742074656D7075;
        inPKT[881]      = 80'hC071732061756775652E;
        inPKT[882]      = 80'hC072204E756C6C612066;
        inPKT[883]      = 80'hC07372696E67696C6C61;
        inPKT[884]      = 80'hC07420656C656966656E;
        inPKT[885]      = 80'hC0756420697073756D20;
        inPKT[886]      = 80'hC0767669766572726120;
        inPKT[887]      = 80'hC0776375727375732E20;
        inPKT[888]      = 80'hC078416C697175616D20;
        inPKT[889]      = 80'hC0796D6178696D757320;
        inPKT[890]      = 80'hC07A6665726D656E7475;
        inPKT[891]      = 80'hC07B6D206E6962682061;
        inPKT[892]      = 80'hC07C6320616363756D73;
        inPKT[893]      = 80'hC07D616E2E204E756C6C;
        inPKT[894]      = 80'hC07E6120666163696C69;
        inPKT[895]      = 80'hC07F73692E2056657374;
        inPKT[896]      = 80'hC0806962756C756D2066;
        inPKT[897]      = 80'hC0816163696C69736973;
        inPKT[898]      = 80'hC082206C656F20656765;
        inPKT[899]      = 80'hC083737461732073656D;
        inPKT[900]      = 80'hC084206D617474697320;
        inPKT[901]      = 80'hC085636F6E6775652E20;
        inPKT[902]      = 80'hC0864D61757269732076;
        inPKT[903]      = 80'hC0876974616520657820;
        inPKT[904]      = 80'hC0886174207269737573;
        inPKT[905]      = 80'hC0892064617069627573;
        inPKT[906]      = 80'hC08A20656C656966656E;
        inPKT[907]      = 80'hC08B642E20496E746567;
        inPKT[908]      = 80'hC08C6572207574206572;
        inPKT[909]      = 80'hC08D6F7320636F6E6775;
        inPKT[910]      = 80'hC08E652C20706F727474;
        inPKT[911]      = 80'hC08F69746F7220616E74;
        inPKT[912]      = 80'hC09065206E6F6E2C2069;
        inPKT[913]      = 80'hC0916E74657264756D20;
        inPKT[914]      = 80'hC092646F6C6F722E0D0A;
        inPKT[915]      = 80'hC0930D0A566573746962;
        inPKT[916]      = 80'hC094756C756D20656C65;
        inPKT[917]      = 80'hC0956966656E64206D61;
        inPKT[918]      = 80'hC0967572697320657520;
        inPKT[919]      = 80'hC0976E69736920646963;
        inPKT[920]      = 80'hC09874756D2067726176;
        inPKT[921]      = 80'hC0996964612E20447569;
        inPKT[922]      = 80'hC09A73206D6F6C6C6973;
        inPKT[923]      = 80'hC09B206469616D207665;
        inPKT[924]      = 80'hC09C6C20656E696D2074;
        inPKT[925]      = 80'hC09D656D7075732C2076;
        inPKT[926]      = 80'hC09E6974616520646170;
        inPKT[927]      = 80'hC09F69627573206D6173;
        inPKT[928]      = 80'hC0A07361207361676974;
        inPKT[929]      = 80'hC0A17469732E204E756C;
        inPKT[930]      = 80'hC0A26C61207574206175;
        inPKT[931]      = 80'hC0A363746F7220746F72;
        inPKT[932]      = 80'hC0A4746F722E204D6F72;
        inPKT[933]      = 80'hC0A5626920736564206C;
        inPKT[934]      = 80'hC0A66F72656D2075726E;
        inPKT[935]      = 80'hC0A7612E204675736365;
        inPKT[936]      = 80'hC0A8206D61747469732C;
        inPKT[937]      = 80'hC0A9206D61676E612061;
        inPKT[938]      = 80'hC0AA6320636F6E64696D;
        inPKT[939]      = 80'hC0AB656E74756D206665;
        inPKT[940]      = 80'hC0AC75676961742C206D;
        inPKT[941]      = 80'hC0AD6173736120647569;
        inPKT[942]      = 80'hC0AE206D6178696D7573;
        inPKT[943]      = 80'hC0AF206E756C6C612C20;
        inPKT[944]      = 80'hC0B0657520616C697175;
        inPKT[945]      = 80'hC0B16574206E65717565;
        inPKT[946]      = 80'hC0B2206D617572697320;
        inPKT[947]      = 80'hC0B36120657261742E20;
        inPKT[948]      = 80'hC0B45175697371756520;
        inPKT[949]      = 80'hC0B5617563746F722065;
        inPKT[950]      = 80'hC0B6737420757420696E;
        inPKT[951]      = 80'hC0B774657264756D2063;
        inPKT[952]      = 80'hC0B86F6E736563746574;
        inPKT[953]      = 80'hC0B975722E20446F6E65;
        inPKT[954]      = 80'hC0BA6320656765742064;
        inPKT[955]      = 80'hC0BB69676E697373696D;
        inPKT[956]      = 80'hC0BC20746F72746F722C;
        inPKT[957]      = 80'hC0BD2068656E64726572;
        inPKT[958]      = 80'hC0BE6974206D61747469;
        inPKT[959]      = 80'hC0BF7320657261742E20;
        inPKT[960]      = 80'hC0C050656C6C656E7465;
        inPKT[961]      = 80'hC0C17371756520686162;
        inPKT[962]      = 80'hC0C26974616E74206D6F;
        inPKT[963]      = 80'hC0C37262692074726973;
        inPKT[964]      = 80'hC0C47469717565207365;
        inPKT[965]      = 80'hC0C56E65637475732065;
        inPKT[966]      = 80'hC0C674206E6574757320;
        inPKT[967]      = 80'hC0C76574206D616C6573;
        inPKT[968]      = 80'hC0C8756164612066616D;
        inPKT[969]      = 80'hC0C96573206163207475;
        inPKT[970]      = 80'hC0CA7270697320656765;
        inPKT[971]      = 80'hC0CB737461732E205175;
        inPKT[972]      = 80'hC0CC6973717565206F72;
        inPKT[973]      = 80'hC0CD6E61726520766172;
        inPKT[974]      = 80'hC0CE6975732074656D70;
        inPKT[975]      = 80'hC0CF75732E0D0A0D0A4D;
        inPKT[976]      = 80'hC0D06F72626920727574;
        inPKT[977]      = 80'hC0D172756D20616E7465;
        inPKT[978]      = 80'hC0D2206E6962682C2061;
        inPKT[979]      = 80'hC0D32076697665727261;
        inPKT[980]      = 80'hC0D4206E756C6C612068;
        inPKT[981]      = 80'hC0D5656E647265726974;
        inPKT[982]      = 80'hC0D620696E2E2050726F;
        inPKT[983]      = 80'hC0D7696E207375736369;
        inPKT[984]      = 80'hC0D87069742065676573;
        inPKT[985]      = 80'hC0D97461732065726174;
        inPKT[986]      = 80'hC0DA2C20757420617563;
        inPKT[987]      = 80'hC0DB746F72206F726369;
        inPKT[988]      = 80'hC0DC206D617474697320;
        inPKT[989]      = 80'hC0DD612E2050656C6C65;
        inPKT[990]      = 80'hC0DE6E74657371756520;
        inPKT[991]      = 80'hC0DF6C75637475732066;
        inPKT[992]      = 80'hC0E072696E67696C6C61;
        inPKT[993]      = 80'hC0E120656C6974207574;
        inPKT[994]      = 80'hC0E2206C6163696E6961;
        inPKT[995]      = 80'hC0E32E20557420657420;
        inPKT[996]      = 80'hC0E46D61737361206E75;
        inPKT[997]      = 80'hC0E56C6C612E20536564;
        inPKT[998]      = 80'hC0E6206174206672696E;
        inPKT[999]      = 80'hC0E767696C6C61206C6F;
        inPKT[1000]     = 80'hC0E872656D2E2050726F;
        inPKT[1001]     = 80'hC0E9696E206772617669;
        inPKT[1002]     = 80'hC0EA646120616363756D;
        inPKT[1003]     = 80'hC0EB73616E2072697375;
        inPKT[1004]     = 80'hC0EC7320736564206269;
        inPKT[1005]     = 80'hC0ED62656E64756D2E20;
        inPKT[1006]     = 80'hC0EE4D616563656E6173;
        inPKT[1007]     = 80'hC0EF206D616C65737561;
        inPKT[1008]     = 80'hC0F06461206F64696F20;
        inPKT[1009]     = 80'hC0F175742076656C6974;
        inPKT[1010]     = 80'hC0F220657569736D6F64;
        inPKT[1011]     = 80'hC0F32064617069627573;
        inPKT[1012]     = 80'hC0F42E0D0A0D0A457469;
        inPKT[1013]     = 80'hC0F5616D20636F6E6775;
        inPKT[1014]     = 80'hC0F665206D6174746973;
        inPKT[1015]     = 80'hC0F720696163756C6973;
        inPKT[1016]     = 80'hC0F82E204D6175726973;
        inPKT[1017]     = 80'hC0F92076697461652065;
        inPKT[1018]     = 80'hC0FA6666696369747572;
        inPKT[1019]     = 80'hC0FB2073656D2E205365;
        inPKT[1020]     = 80'hC0FC642070756C76696E;
        inPKT[1021]     = 80'hC0FD617220646F6C6F72;
        inPKT[1022]     = 80'hC0FE207574206D692065;
        inPKT[1023]     = 80'hC0FF7569736D6F642068;
        inPKT[1024]     = 80'hC000656E647265726974;
        inPKT[1025]     = 80'hC0012E204E756C6C616D;
        inPKT[1026]     = 80'hC0022061742067726176;
        inPKT[1027]     = 80'hC00369646120646F6C6F;
        inPKT[1028]     = 80'hC004722E204D6F726269;
        inPKT[1029]     = 80'hC005206C656F20747572;
        inPKT[1030]     = 80'hC0067069732C20636F6E;
        inPKT[1031]     = 80'hC007677565206E656320;
        inPKT[1032]     = 80'hC008616C697175616D20;
        inPKT[1033]     = 80'hC00975742C20636F6D6D;
        inPKT[1034]     = 80'hC00A6F646F20696E206E;
        inPKT[1035]     = 80'hC00B756E632E204E756C;
        inPKT[1036]     = 80'hC00C6C61206174206661;
        inPKT[1037]     = 80'hC00D756369627573206C;
        inPKT[1038]     = 80'hC00E656F2C2065752066;
        inPKT[1039]     = 80'hC00F657567696174206C;
        inPKT[1040]     = 80'hC010616375732E204675;
        inPKT[1041]     = 80'hC011736365206E6F6E20;
        inPKT[1042]     = 80'hC0126567657374617320;
        inPKT[1043]     = 80'hC0137475727069732E20;
        inPKT[1044]     = 80'hC0145175697371756520;
        inPKT[1045]     = 80'hC0157669746165206970;
        inPKT[1046]     = 80'hC01673756D206D692E20;
        inPKT[1047]     = 80'hC0174E756E63206E6F6E;
        inPKT[1048]     = 80'hC018206F726369207369;
        inPKT[1049]     = 80'hC0197420616D6574206E;
        inPKT[1050]     = 80'hC01A6973692076617269;
        inPKT[1051]     = 80'hC01B757320706F727474;
        inPKT[1052]     = 80'hC01C69746F7220696E20;
        inPKT[1053]     = 80'hC01D76756C7075746174;
        inPKT[1054]     = 80'hC01E6520746F72746F72;
        inPKT[1055]     = 80'hC01F2E204E756E632063;
        inPKT[1056]     = 80'hC0206F6E76616C6C6973;
        inPKT[1057]     = 80'hC0212067726176696461;
        inPKT[1058]     = 80'hC022206469616D206120;
        inPKT[1059]     = 80'hC023756C747269636965;
        inPKT[1060]     = 80'hC024732E205175697371;
        inPKT[1061]     = 80'hC0257565206575206A75;
        inPKT[1062]     = 80'hC02673746F20636F6E64;
        inPKT[1063]     = 80'hC027696D656E74756D2C;
        inPKT[1064]     = 80'hC0282076617269757320;
        inPKT[1065]     = 80'hC0296469616D2076656C;
        inPKT[1066]     = 80'hC02A2C20766573746962;
        inPKT[1067]     = 80'hC02B756C756D206D6173;
        inPKT[1068]     = 80'hC02C73612E0D0A0D0A50;
        inPKT[1069]     = 80'hC02D656C6C656E746573;
        inPKT[1070]     = 80'hC02E7175652070656C6C;
        inPKT[1071]     = 80'hC02F656E746573717565;
        inPKT[1072]     = 80'hC0302073617069656E20;
        inPKT[1073]     = 80'hC0316E657175652C2061;
        inPKT[1074]     = 80'hC0327563746F72206D61;
        inPKT[1075]     = 80'hC0336C65737561646120;
        inPKT[1076]     = 80'hC034657261742068656E;
        inPKT[1077]     = 80'hC035647265726974206E;
        inPKT[1078]     = 80'hC03665632E204E756C6C;
        inPKT[1079]     = 80'hC0376120706C61636572;
        inPKT[1080]     = 80'hC0386174206469616D20;
        inPKT[1081]     = 80'hC03968656E6472657269;
        inPKT[1082]     = 80'hC03A74206D6173736120;
        inPKT[1083]     = 80'hC03B626962656E64756D;
        inPKT[1084]     = 80'hC03C2C2061206D6F6C65;
        inPKT[1085]     = 80'hC03D737469652066656C;
        inPKT[1086]     = 80'hC03E69732068656E6472;
        inPKT[1087]     = 80'hC03F657269742E204D61;
        inPKT[1088]     = 80'hC0407572697320657569;
        inPKT[1089]     = 80'hC041736D6F642076656E;
        inPKT[1090]     = 80'hC042656E61746973206A;
        inPKT[1091]     = 80'hC0437573746F2C207574;
        inPKT[1092]     = 80'hC04420617563746F7220;
        inPKT[1093]     = 80'hC045656C697420616C69;
        inPKT[1094]     = 80'hC046717565742075742E;
        inPKT[1095]     = 80'hC0472046757363652061;
        inPKT[1096]     = 80'hC0486C69717565742C20;
        inPKT[1097]     = 80'hC0497175616D20757420;
        inPKT[1098]     = 80'hC04A6469676E69737369;
        inPKT[1099]     = 80'hC04B6D2068656E647265;
        inPKT[1100]     = 80'hC04C7269742C206D6175;
        inPKT[1101]     = 80'hC04D7269732074757270;
        inPKT[1102]     = 80'hC04E6973206469676E69;
        inPKT[1103]     = 80'hC04F7373696D20746F72;
        inPKT[1104]     = 80'hC050746F722C20656765;
        inPKT[1105]     = 80'hC051742070656C6C656E;
        inPKT[1106]     = 80'hC0527465737175652076;
        inPKT[1107]     = 80'hC053656C6974206F7263;
        inPKT[1108]     = 80'hC05469206E6563207175;
        inPKT[1109]     = 80'hC055616D2E204E756E63;
        inPKT[1110]     = 80'hC0562065676573746173;
        inPKT[1111]     = 80'hC0572070656C6C656E74;
        inPKT[1112]     = 80'hC0586573717565207269;
        inPKT[1113]     = 80'hC0597375732E20437572;
        inPKT[1114]     = 80'hC05A6162697475722073;
        inPKT[1115]     = 80'hC05B7573636970697420;
        inPKT[1116]     = 80'hC05C74656D707573206C;
        inPKT[1117]     = 80'hC05D616375732C206567;
        inPKT[1118]     = 80'hC05E6574207072657469;
        inPKT[1119]     = 80'hC05F756D20656C697420;
        inPKT[1120]     = 80'hC06074696E636964756E;
        inPKT[1121]     = 80'hC06174206E6F6E2E2043;
        inPKT[1122]     = 80'hC0627261732075726E61;
        inPKT[1123]     = 80'hC063206C6F72656D2C20;
        inPKT[1124]     = 80'hC064706C616365726174;
        inPKT[1125]     = 80'hC06520766F6C75747061;
        inPKT[1126]     = 80'hC0667420696D70657264;
        inPKT[1127]     = 80'hC0676965742073697420;
        inPKT[1128]     = 80'hC068616D65742C206567;
        inPKT[1129]     = 80'hC0696573746173207665;
        inPKT[1130]     = 80'hC06A6C206F7263692E0D;
        inPKT[1131]     = 80'hC06B0A0D0A50656C6C65;
        inPKT[1132]     = 80'hC06C6E74657371756520;
        inPKT[1133]     = 80'hC06D736F64616C657320;
        inPKT[1134]     = 80'hC06E6665726D656E7475;
        inPKT[1135]     = 80'hC06F6D206E69736C2C20;
        inPKT[1136]     = 80'hC0706174206672696E67;
        inPKT[1137]     = 80'hC071696C6C6120647569;
        inPKT[1138]     = 80'hC0722073656D70657220;
        inPKT[1139]     = 80'hC0736665726D656E7475;
        inPKT[1140]     = 80'hC0746D2E204E756C6C61;
        inPKT[1141]     = 80'hC0756D20706C61636572;
        inPKT[1142]     = 80'hC07661742076656C206D;
        inPKT[1143]     = 80'hC077692068656E647265;
        inPKT[1144]     = 80'hC07872697420656C656D;
        inPKT[1145]     = 80'hC079656E74756D2E2045;
        inPKT[1146]     = 80'hC07A7469616D206E6F6E;
        inPKT[1147]     = 80'hC07B20697073756D2065;
        inPKT[1148]     = 80'hC07C782E204E616D2061;
        inPKT[1149]     = 80'hC07D63207363656C6572;
        inPKT[1150]     = 80'hC07E6973717565206E69;
        inPKT[1151]     = 80'hC07F62682C2076656C20;
        inPKT[1152]     = 80'hC080666163696C697369;
        inPKT[1153]     = 80'hC08173206D692E20446F;
        inPKT[1154]     = 80'hC0826E65632065676573;
        inPKT[1155]     = 80'hC083746173206C616F72;
        inPKT[1156]     = 80'hC0846565742065726F73;
        inPKT[1157]     = 80'hC0852C20656765742076;
        inPKT[1158]     = 80'hC0866F6C757470617420;
        inPKT[1159]     = 80'hC0876D657475732E2050;
        inPKT[1160]     = 80'hC08872616573656E7420;
        inPKT[1161]     = 80'hC089616363756D73616E;
        inPKT[1162]     = 80'hC08A20626962656E6475;
        inPKT[1163]     = 80'hC08B6D206E69736C206E;
        inPKT[1164]     = 80'hC08C65632076656E656E;
        inPKT[1165]     = 80'hC08D617469732E205365;
        inPKT[1166]     = 80'hC08E642072757472756D;
        inPKT[1167]     = 80'hC08F206D692061207375;
        inPKT[1168]     = 80'hC0907363697069742070;
        inPKT[1169]     = 80'hC091686172657472612E;
        inPKT[1170]     = 80'hC0922053656420736974;
        inPKT[1171]     = 80'hC09320616D657420696E;
        inPKT[1172]     = 80'hC09474657264756D2074;
        inPKT[1173]     = 80'hC09575727069732E2041;
        inPKT[1174]     = 80'hC0966C697175616D2065;
        inPKT[1175]     = 80'hC09775206E6962682074;
        inPKT[1176]     = 80'hC0986F72746F722E2044;
        inPKT[1177]     = 80'hC0996F6E656320666175;
        inPKT[1178]     = 80'hC09A6369627573206461;
        inPKT[1179]     = 80'hC09B7069627573206E69;
        inPKT[1180]     = 80'hC09C73692C2073656420;
        inPKT[1181]     = 80'hC09D6C616F7265657420;
        inPKT[1182]     = 80'hC09E6F72636920736365;
        inPKT[1183]     = 80'hC09F6C65726973717565;
        inPKT[1184]     = 80'hC0A020696E2E0D0A0D0A;
        inPKT[1185]     = 80'hC0A14D61757269732069;
        inPKT[1186]     = 80'hC0A26E2066656C697320;
        inPKT[1187]     = 80'hC0A36665726D656E7475;
        inPKT[1188]     = 80'hC0A46D2C20636F6E7661;
        inPKT[1189]     = 80'hC0A56C6C697320617567;
        inPKT[1190]     = 80'hC0A675652076656C2C20;
        inPKT[1191]     = 80'hC0A7706F737565726520;
        inPKT[1192]     = 80'hC0A86D692E2050656C6C;
        inPKT[1193]     = 80'hC0A9656E746573717565;
        inPKT[1194]     = 80'hC0AA207363656C657269;
        inPKT[1195]     = 80'hC0AB737175652072686F;
        inPKT[1196]     = 80'hC0AC6E637573206A7573;
        inPKT[1197]     = 80'hC0AD746F2C2065752070;
        inPKT[1198]     = 80'hC0AE756C76696E617220;
        inPKT[1199]     = 80'hC0AF656E696D2070756C;
        inPKT[1200]     = 80'hC0B076696E6172207665;
        inPKT[1201]     = 80'hC0B16C2E204D61656365;
        inPKT[1202]     = 80'hC0B26E61732070686172;
        inPKT[1203]     = 80'hC0B365747261206C6962;
        inPKT[1204]     = 80'hC0B465726F206D61676E;
        inPKT[1205]     = 80'hC0B5612C20616320736F;
        inPKT[1206]     = 80'hC0B66C6C696369747564;
        inPKT[1207]     = 80'hC0B7696E206C656F206D;
        inPKT[1208]     = 80'hC0B86F6C6C6973206E6F;
        inPKT[1209]     = 80'hC0B96E2E204E756C6C61;
        inPKT[1210]     = 80'hC0BA20656C656D656E74;
        inPKT[1211]     = 80'hC0BB756D206F726E6172;
        inPKT[1212]     = 80'hC0BC6520656765737461;
        inPKT[1213]     = 80'hC0BD732E20436C617373;
        inPKT[1214]     = 80'hC0BE20617074656E7420;
        inPKT[1215]     = 80'hC0BF7461636974692073;
        inPKT[1216]     = 80'hC0C06F63696F73717520;
        inPKT[1217]     = 80'hC0C16164206C69746F72;
        inPKT[1218]     = 80'hC0C26120746F72717565;
        inPKT[1219]     = 80'hC0C36E74207065722063;
        inPKT[1220]     = 80'hC0C46F6E75626961206E;
        inPKT[1221]     = 80'hC0C56F737472612C2070;
        inPKT[1222]     = 80'hC0C6657220696E636570;
        inPKT[1223]     = 80'hC0C7746F732068696D65;
        inPKT[1224]     = 80'hC0C86E61656F732E2050;
        inPKT[1225]     = 80'hC0C972616573656E7420;
        inPKT[1226]     = 80'hC0CA6175677565206D61;
        inPKT[1227]     = 80'hC0CB757269732C207268;
        inPKT[1228]     = 80'hC0CC6F6E637573207175;
        inPKT[1229]     = 80'hC0CD697320657374206E;
        inPKT[1230]     = 80'hC0CE6F6E2C206D6F6C6C;
        inPKT[1231]     = 80'hC0CF697320636F6E7661;
        inPKT[1232]     = 80'hC0D06C6C69732066656C;
        inPKT[1233]     = 80'hC0D169732E2053757370;
        inPKT[1234]     = 80'hC0D2656E646973736520;
        inPKT[1235]     = 80'hC0D3666163696C697369;
        inPKT[1236]     = 80'hC0D4732C206F72636920;
        inPKT[1237]     = 80'hC0D57669746165206C61;
        inPKT[1238]     = 80'hC0D663696E6961207465;
        inPKT[1239]     = 80'hC0D76D706F722C206C65;
        inPKT[1240]     = 80'hC0D86374757320736170;
        inPKT[1241]     = 80'hC0D969656E206D617474;
        inPKT[1242]     = 80'hC0DA6973207269737573;
        inPKT[1243]     = 80'hC0DB2C206E6F6E207361;
        inPKT[1244]     = 80'hC0DC6769747469732065;
        inPKT[1245]     = 80'hC0DD6C6974206E657175;
        inPKT[1246]     = 80'hC0DE652071756973206A;
        inPKT[1247]     = 80'hC0DF7573746F2E20446F;
        inPKT[1248]     = 80'hC0E06E6563206D616C65;
        inPKT[1249]     = 80'hC0E17375616461206C61;
        inPKT[1250]     = 80'hC0E263696E6961206475;
        inPKT[1251]     = 80'hC0E3692E205068617365;
        inPKT[1252]     = 80'hC0E46C6C75732068656E;
        inPKT[1253]     = 80'hC0E5647265726974206D;
        inPKT[1254]     = 80'hC0E66175726973206D61;
        inPKT[1255]     = 80'hC0E7757269732C207365;
        inPKT[1256]     = 80'hC0E864206672696E6769;
        inPKT[1257]     = 80'hC0E96C6C61206C696265;
        inPKT[1258]     = 80'hC0EA726F206672696E67;
        inPKT[1259]     = 80'hC0EB696C6C6120696E2E;
        inPKT[1260]     = 80'hC0EC2053656420617420;
        inPKT[1261]     = 80'hC0ED6C6967756C612069;
        inPKT[1262]     = 80'hC0EE6E206A7573746F20;
        inPKT[1263]     = 80'hC0EF66696E6962757320;
        inPKT[1264]     = 80'hC0F076756C7075746174;
        inPKT[1265]     = 80'hC0F1652E204E756E6320;
        inPKT[1266]     = 80'hC0F2637572737573206E;
        inPKT[1267]     = 80'hC0F36571756520736974;
        inPKT[1268]     = 80'hC0F420616D6574206172;
        inPKT[1269]     = 80'hC0F563752074696E6369;
        inPKT[1270]     = 80'hC0F664756E742C207669;
        inPKT[1271]     = 80'hC0F77461652070686172;
        inPKT[1272]     = 80'hC0F8657472612073656D;
        inPKT[1273]     = 80'hC0F920706F7274746974;
        inPKT[1274]     = 80'hC0FA6F722E20416C6971;
        inPKT[1275]     = 80'hC0FB75616D206D617474;
        inPKT[1276]     = 80'hC0FC69732C206A757374;
        inPKT[1277]     = 80'hC0FD6F206E6F6E206575;
        inPKT[1278]     = 80'hC0FE69736D6F6420636F;
        inPKT[1279]     = 80'hC0FF6E76616C6C69732C;
        inPKT[1280]     = 80'hC000206E756E63206D69;
        inPKT[1281]     = 80'hC00120636F6E73657175;
        inPKT[1282]     = 80'hC0026174206573742C20;
        inPKT[1283]     = 80'hC0036E656320736F6C6C;
        inPKT[1284]     = 80'hC004696369747564696E;
        inPKT[1285]     = 80'hC005206C656374757320;
        inPKT[1286]     = 80'hC00673617069656E2076;
        inPKT[1287]     = 80'hC007656C206F64696F2E;
        inPKT[1288]     = 80'hC00820496E2074656D70;
        inPKT[1289]     = 80'hC0096F72206572617420;
        inPKT[1290]     = 80'hC00A646F6C6F722C2073;
        inPKT[1291]     = 80'hC00B6564207665686963;
        inPKT[1292]     = 80'hC00C756C612075726E61;
        inPKT[1293]     = 80'hC00D20636F6E73657175;
        inPKT[1294]     = 80'hC00E6174207365642E0D;
        inPKT[1295]     = 80'hC00F0A0D0A4E616D2072;
        inPKT[1296]     = 80'hC010686F6E6375732069;
        inPKT[1297]     = 80'hC01164206D6175726973;
        inPKT[1298]     = 80'hC012206E656320646967;
        inPKT[1299]     = 80'hC0136E697373696D2E20;
        inPKT[1300]     = 80'hC014496E20696D706572;
        inPKT[1301]     = 80'hC0156469657420756C74;
        inPKT[1302]     = 80'hC0167269636573206572;
        inPKT[1303]     = 80'hC0176174206E65632073;
        inPKT[1304]     = 80'hC0186F6C6C6963697475;
        inPKT[1305]     = 80'hC01964696E2E20496E74;
        inPKT[1306]     = 80'hC01A6567657220736564;
        inPKT[1307]     = 80'hC01B20636F6E64696D65;
        inPKT[1308]     = 80'hC01C6E74756D2065726F;
        inPKT[1309]     = 80'hC01D732E20446F6E6563;
        inPKT[1310]     = 80'hC01E2065676574206E75;
        inPKT[1311]     = 80'hC01F6E63206964206D61;
        inPKT[1312]     = 80'hC0207572697320747269;
        inPKT[1313]     = 80'hC0217374697175652070;
        inPKT[1314]     = 80'hC0226F72747469746F72;
        inPKT[1315]     = 80'hC023206C616F72656574;
        inPKT[1316]     = 80'hC024207669746165206D;
        inPKT[1317]     = 80'hC025657475732E204E75;
        inPKT[1318]     = 80'hC0266C6C612066616369;
        inPKT[1319]     = 80'hC0276C6973692E204E75;
        inPKT[1320]     = 80'hC0286C6C616D20657520;
        inPKT[1321]     = 80'hC0296C61637573206120;
        inPKT[1322]     = 80'hC02A6469616D20747269;
        inPKT[1323]     = 80'hC02B7374697175652065;
        inPKT[1324]     = 80'hC02C676573746173206E;
        inPKT[1325]     = 80'hC02D6F6E20696163756C;
        inPKT[1326]     = 80'hC02E6973206D65747573;
        inPKT[1327]     = 80'hC02F2E20416C69717561;
        inPKT[1328]     = 80'hC0306D20696E2074656D;
        inPKT[1329]     = 80'hC031706F722065726174;
        inPKT[1330]     = 80'hC0322C20696420636F6E;
        inPKT[1331]     = 80'hC033677565206D617373;
        inPKT[1332]     = 80'hC034612E20566976616D;
        inPKT[1333]     = 80'hC03575732076656C2074;
        inPKT[1334]     = 80'hC0366F72746F72207669;
        inPKT[1335]     = 80'hC037746165206E696268;
        inPKT[1336]     = 80'hC03820636F6D6D6F646F;
        inPKT[1337]     = 80'hC039206C6F626F727469;
        inPKT[1338]     = 80'hC03A7320717569732061;
        inPKT[1339]     = 80'hC03B20697073756D2E20;
        inPKT[1340]     = 80'hC03C50726F696E20766F;
        inPKT[1341]     = 80'hC03D6C75747061742071;
        inPKT[1342]     = 80'hC03E75616D206E6F6E20;
        inPKT[1343]     = 80'hC03F66656C6973207465;
        inPKT[1344]     = 80'hC0406D7075732C206964;
        inPKT[1345]     = 80'hC04120706F7375657265;
        inPKT[1346]     = 80'hC04220646F6C6F722074;
        inPKT[1347]     = 80'hC043656D706F722E2050;
        inPKT[1348]     = 80'hC04472616573656E7420;
        inPKT[1349]     = 80'hC0457669746165207469;
        inPKT[1350]     = 80'hC0466E636964756E7420;
        inPKT[1351]     = 80'hC04773617069656E2E20;
        inPKT[1352]     = 80'hC0484D616563656E6173;
        inPKT[1353]     = 80'hC04920666163696C6973;
        inPKT[1354]     = 80'hC04A6973206D61747469;
        inPKT[1355]     = 80'hC04B7320616E74652071;
        inPKT[1356]     = 80'hC04C7569732076617269;
        inPKT[1357]     = 80'hC04D75732E20446F6E65;
        inPKT[1358]     = 80'hC04E632070656C6C656E;
        inPKT[1359]     = 80'hC04F7465737175652065;
        inPKT[1360]     = 80'hC050726F732066657567;
        inPKT[1361]     = 80'hC0516961742074696E63;
        inPKT[1362]     = 80'hC0526964756E7420636F;
        inPKT[1363]     = 80'hC0536E64696D656E7475;
        inPKT[1364]     = 80'hC0546D2E2050726F696E;
        inPKT[1365]     = 80'hC0552066617563696275;
        inPKT[1366]     = 80'hC0567320766F6C757470;
        inPKT[1367]     = 80'hC0576174206D69207365;
        inPKT[1368]     = 80'hC0586420736167697474;
        inPKT[1369]     = 80'hC05969732E0D0A0D0A44;
        inPKT[1370]     = 80'hC05A7569732067726176;
        inPKT[1371]     = 80'hC05B69646120656C656D;
        inPKT[1372]     = 80'hC05C656E74756D20696E;
        inPKT[1373]     = 80'hC05D74657264756D2E20;
        inPKT[1374]     = 80'hC05E50726F696E207369;
        inPKT[1375]     = 80'hC05F7420616D65742071;
        inPKT[1376]     = 80'hC06075616D206C696775;
        inPKT[1377]     = 80'hC0616C612E2050686173;
        inPKT[1378]     = 80'hC062656C6C757320636F;
        inPKT[1379]     = 80'hC0636D6D6F646F2C2075;
        inPKT[1380]     = 80'hC064726E6120696E2063;
        inPKT[1381]     = 80'hC0656F6E67756520766F;
        inPKT[1382]     = 80'hC0666C75747061742C20;
        inPKT[1383]     = 80'hC0676C6967756C612065;
        inPKT[1384]     = 80'hC0687820706861726574;
        inPKT[1385]     = 80'hC0697261206C6967756C;
        inPKT[1386]     = 80'hC06A612C20696E206469;
        inPKT[1387]     = 80'hC06B6374756D206D6167;
        inPKT[1388]     = 80'hC06C6E61206F72636920;
        inPKT[1389]     = 80'hC06D6E6563206D617572;
        inPKT[1390]     = 80'hC06E69732E204E756E63;
        inPKT[1391]     = 80'hC06F20617563746F7220;
        inPKT[1392]     = 80'hC070636F6E7365637465;
        inPKT[1393]     = 80'hC07174757220766F6C75;
        inPKT[1394]     = 80'hC072747061742E204D6F;
        inPKT[1395]     = 80'hC0737262692074696E63;
        inPKT[1396]     = 80'hC0746964756E74206E69;
        inPKT[1397]     = 80'hC075626820757420656E;
        inPKT[1398]     = 80'hC076696D206566666963;
        inPKT[1399]     = 80'hC0776974757220677261;
        inPKT[1400]     = 80'hC078766964612E204375;
        inPKT[1401]     = 80'hC0797261626974757220;
        inPKT[1402]     = 80'hC07A7669746165207175;
        inPKT[1403]     = 80'hC07B616D2065726F732E;
        inPKT[1404]     = 80'hC07C2044756973206672;
        inPKT[1405]     = 80'hC07D696E67696C6C6120;
        inPKT[1406]     = 80'hC07E616320746F72746F;
        inPKT[1407]     = 80'hC07F7220696E2074696E;
        inPKT[1408]     = 80'hC080636964756E742E20;
        inPKT[1409]     = 80'hC0814E756E632076656C;
        inPKT[1410]     = 80'hC082206D617572697320;
        inPKT[1411]     = 80'hC08372697375732E2044;
        inPKT[1412]     = 80'hC0846F6E656320656C65;
        inPKT[1413]     = 80'hC0856966656E64206C69;
        inPKT[1414]     = 80'hC08667756C6120736167;
        inPKT[1415]     = 80'hC0876974746973206E69;
        inPKT[1416]     = 80'hC08873692066696E6962;
        inPKT[1417]     = 80'hC08975732C2061207363;
        inPKT[1418]     = 80'hC08A656C657269737175;
        inPKT[1419]     = 80'hC08B65206C696265726F;
        inPKT[1420]     = 80'hC08C2070656C6C656E74;
        inPKT[1421]     = 80'hC08D65737175652E2056;
        inPKT[1422]     = 80'hC08E6573746962756C75;
        inPKT[1423]     = 80'hC08F6D20747269737469;
        inPKT[1424]     = 80'hC090717565206D617373;
        inPKT[1425]     = 80'hC09161206E6962682C20;
        inPKT[1426]     = 80'hC0926174207665737469;
        inPKT[1427]     = 80'hC09362756C756D206D61;
        inPKT[1428]     = 80'hC094676E612066696E69;
        inPKT[1429]     = 80'hC0956275732065752E0D;
        inPKT[1430]     = 80'hC0960A0D0A4375726162;
        inPKT[1431]     = 80'hC0976974757220696D70;
        inPKT[1432]     = 80'hC0986572646965742070;
        inPKT[1433]     = 80'hC0997572757320656765;
        inPKT[1434]     = 80'hC09A74206E756E632075;
        inPKT[1435]     = 80'hC09B6C7472696365732C;
        inPKT[1436]     = 80'hC09C2076697461652076;
        inPKT[1437]     = 80'hC09D656E656E61746973;
        inPKT[1438]     = 80'hC09E206D617373612063;
        inPKT[1439]     = 80'hC09F6F6D6D6F646F2E20;
        inPKT[1440]     = 80'hC0A050656C6C656E7465;
        inPKT[1441]     = 80'hC0A17371756520686162;
        inPKT[1442]     = 80'hC0A26974616E74206D6F;
        inPKT[1443]     = 80'hC0A37262692074726973;
        inPKT[1444]     = 80'hC0A47469717565207365;
        inPKT[1445]     = 80'hC0A56E65637475732065;
        inPKT[1446]     = 80'hC0A674206E6574757320;
        inPKT[1447]     = 80'hC0A76574206D616C6573;
        inPKT[1448]     = 80'hC0A8756164612066616D;
        inPKT[1449]     = 80'hC0A96573206163207475;
        inPKT[1450]     = 80'hC0AA7270697320656765;
        inPKT[1451]     = 80'hC0AB737461732E20496E;
        inPKT[1452]     = 80'hC0AC206665726D656E74;
        inPKT[1453]     = 80'hC0AD756D206174207572;
        inPKT[1454]     = 80'hC0AE6E61206E6F6E2063;
        inPKT[1455]     = 80'hC0AF6F6E76616C6C6973;
        inPKT[1456]     = 80'hC0B02E20446F6E656320;
        inPKT[1457]     = 80'hC0B16163206175677565;
        inPKT[1458]     = 80'hC0B2206A7573746F2E20;
        inPKT[1459]     = 80'hC0B3496E20617420656C;
        inPKT[1460]     = 80'hC0B46974206574206172;
        inPKT[1461]     = 80'hC0B56375206D6178696D;
        inPKT[1462]     = 80'hC0B67573206C75637475;
        inPKT[1463]     = 80'hC0B7732E204675736365;
        inPKT[1464]     = 80'hC0B820657569736D6F64;
        inPKT[1465]     = 80'hC0B9206E756E63206E65;
        inPKT[1466]     = 80'hC0BA632076656E656E61;
        inPKT[1467]     = 80'hC0BB7469732061756374;
        inPKT[1468]     = 80'hC0BC6F722E204C6F7265;
        inPKT[1469]     = 80'hC0BD6D20697073756D20;
        inPKT[1470]     = 80'hC0BE646F6C6F72207369;
        inPKT[1471]     = 80'hC0BF7420616D65742C20;
        inPKT[1472]     = 80'hC0C0636F6E7365637465;
        inPKT[1473]     = 80'hC0C17475722061646970;
        inPKT[1474]     = 80'hC0C2697363696E672065;
        inPKT[1475]     = 80'hC0C36C69742E20446F6E;
        inPKT[1476]     = 80'hC0C46563206469637475;
        inPKT[1477]     = 80'hC0C56D2074656D706F72;
        inPKT[1478]     = 80'hC0C62072757472756D2E;
        inPKT[1479]     = 80'hC0C72053656420656C65;
        inPKT[1480]     = 80'hC0C86966656E64206469;
        inPKT[1481]     = 80'hC0C9616D206964206D61;
        inPKT[1482]     = 80'hC0CA73736120696D7065;
        inPKT[1483]     = 80'hC0CB72646965742C2061;
        inPKT[1484]     = 80'hC0CC63206F726E617265;
        inPKT[1485]     = 80'hC0CD206C696265726F20;
        inPKT[1486]     = 80'hC0CE656C656966656E64;
        inPKT[1487]     = 80'hC0CF2E204D616563656E;
        inPKT[1488]     = 80'hC0D06173206F726E6172;
        inPKT[1489]     = 80'hC0D165206D6574757320;
        inPKT[1490]     = 80'hC0D26E756C6C612C2073;
        inPKT[1491]     = 80'hC0D3697420616D657420;
        inPKT[1492]     = 80'hC0D46665726D656E7475;
        inPKT[1493]     = 80'hC0D56D20656C69742061;
        inPKT[1494]     = 80'hC0D66C697175616D2069;
        inPKT[1495]     = 80'hC0D7642E20446F6E6563;
        inPKT[1496]     = 80'hC0D820756C7472696365;
        inPKT[1497]     = 80'hC0D97320746F72746F72;
        inPKT[1498]     = 80'hC0DA20617420616E7465;
        inPKT[1499]     = 80'hC0DB2068656E64726572;
        inPKT[1500]     = 80'hC0DC69742C2065752073;
        inPKT[1501]     = 80'hC0DD6167697474697320;
        inPKT[1502]     = 80'hC0DE6A7573746F20756C;
        inPKT[1503]     = 80'hC0DF7472696365732E0D;
        inPKT[1504]     = 80'hC0E00A0D0A5072616573;
        inPKT[1505]     = 80'hC0E1656E74206C756374;
        inPKT[1506]     = 80'hC0E27573207072657469;
        inPKT[1507]     = 80'hC0E3756D206E65717565;
        inPKT[1508]     = 80'hC0E42C2073697420616D;
        inPKT[1509]     = 80'hC0E565742070656C6C65;
        inPKT[1510]     = 80'hC0E66E74657371756520;
        inPKT[1511]     = 80'hC0E76D61757269732065;
        inPKT[1512]     = 80'hC0E86C656D656E74756D;
        inPKT[1513]     = 80'hC0E9206E6F6E2E205574;
        inPKT[1514]     = 80'hC0EA20626C616E646974;
        inPKT[1515]     = 80'hC0EB2070686172657472;
        inPKT[1516]     = 80'hC0EC61206F64696F206E;
        inPKT[1517]     = 80'hC0ED6F6E20657569736D;
        inPKT[1518]     = 80'hC0EE6F642E2051756973;
        inPKT[1519]     = 80'hC0EF7175652076697461;
        inPKT[1520]     = 80'hC0F065206C656F20616C;
        inPKT[1521]     = 80'hC0F1697175616D2C2073;
        inPKT[1522]     = 80'hC0F26F64616C65732074;
        inPKT[1523]     = 80'hC0F3656C6C7573206964;
        inPKT[1524]     = 80'hC0F42C20696163756C69;
        inPKT[1525]     = 80'hC0F573206D6175726973;
        inPKT[1526]     = 80'hC0F62E204E616D206566;
        inPKT[1527]     = 80'hC0F76669636974757220;
        inPKT[1528]     = 80'hC0F8696E207075727573;
        inPKT[1529]     = 80'hC0F92073656420616363;
        inPKT[1530]     = 80'hC0FA756D73616E2E204D;
        inPKT[1531]     = 80'hC0FB616563656E617320;
        inPKT[1532]     = 80'hC0FC73697420616D6574;
        inPKT[1533]     = 80'hC0FD2063757273757320;
        inPKT[1534]     = 80'hC0FE66656C69732E2051;
        inPKT[1535]     = 80'hC0FF7569737175652066;
        inPKT[1536]     = 80'hC000617563696275732C;
        inPKT[1537]     = 80'hC0012064756920657420;
        inPKT[1538]     = 80'hC002617563746F72206C;
        inPKT[1539]     = 80'hC00375637475732C2061;
        inPKT[1540]     = 80'hC0046E74652065726174;
        inPKT[1541]     = 80'hC00520706F7375657265;
        inPKT[1542]     = 80'hC0062065726F732C2075;
        inPKT[1543]     = 80'hC0077420636F6E76616C;
        inPKT[1544]     = 80'hC0086C6973206D657475;
        inPKT[1545]     = 80'hC00973206C6563747573;
        inPKT[1546]     = 80'hC00A207669746165206C;
        inPKT[1547]     = 80'hC00B656F2E2053757370;
        inPKT[1548]     = 80'hC00C656E646973736520;
        inPKT[1549]     = 80'hC00D706F74656E74692E;
        inPKT[1550]     = 80'hC00E2043726173206574;
        inPKT[1551]     = 80'hC00F20646F6C6F72206E;
        inPKT[1552]     = 80'hC0106F6E2075726E6120;
        inPKT[1553]     = 80'hC0117363656C65726973;
        inPKT[1554]     = 80'hC0127175652074726973;
        inPKT[1555]     = 80'hC01374697175652E2043;
        inPKT[1556]     = 80'hC0147261732072757472;
        inPKT[1557]     = 80'hC015756D206E65632076;
        inPKT[1558]     = 80'hC016656C697420616320;
        inPKT[1559]     = 80'hC0177361676974746973;
        inPKT[1560]     = 80'hC0182E20446F6E656320;
        inPKT[1561]     = 80'hC019656C656966656E64;
        inPKT[1562]     = 80'hC01A2C206C6163757320;
        inPKT[1563]     = 80'hC01B7365642067726176;
        inPKT[1564]     = 80'hC01C696461206D616C65;
        inPKT[1565]     = 80'hC01D73756164612C2065;
        inPKT[1566]     = 80'hC01E7820616E74652070;
        inPKT[1567]     = 80'hC01F6C61636572617420;
        inPKT[1568]     = 80'hC0206C65637475732C20;
        inPKT[1569]     = 80'hC0216567657420636F6E;
        inPKT[1570]     = 80'hC022677565206D617373;
        inPKT[1571]     = 80'hC02361206D6574757320;
        inPKT[1572]     = 80'hC0246964206C61637573;
        inPKT[1573]     = 80'hC0252E2053757370656E;
        inPKT[1574]     = 80'hC0266469737365206964;
        inPKT[1575]     = 80'hC0272072757472756D20;
        inPKT[1576]     = 80'hC0286C65637475732E20;
        inPKT[1577]     = 80'hC0294675736365206D61;
        inPKT[1578]     = 80'hC02A78696D7573207365;
        inPKT[1579]     = 80'hC02B64206C6967756C61;
        inPKT[1580]     = 80'hC02C2073656420766976;
        inPKT[1581]     = 80'hC02D657272612E204E61;
        inPKT[1582]     = 80'hC02E6D206C7563747573;
        inPKT[1583]     = 80'hC02F206469616D20616E;
        inPKT[1584]     = 80'hC03074652C2076697461;
        inPKT[1585]     = 80'hC03165206F726E617265;
        inPKT[1586]     = 80'hC032206E657175652076;
        inPKT[1587]     = 80'hC0336172697573206567;
        inPKT[1588]     = 80'hC03465742E0D0A0D0A50;
        inPKT[1589]     = 80'hC035656C6C656E746573;
        inPKT[1590]     = 80'hC0367175652061742065;
        inPKT[1591]     = 80'hC0376C6974206E696268;
        inPKT[1592]     = 80'hC0382E20566573746962;
        inPKT[1593]     = 80'hC039756C756D20616E74;
        inPKT[1594]     = 80'hC03A6520697073756D20;
        inPKT[1595]     = 80'hC03B7072696D69732069;
        inPKT[1596]     = 80'hC03C6E20666175636962;
        inPKT[1597]     = 80'hC03D7573206F72636920;
        inPKT[1598]     = 80'hC03E6C75637475732065;
        inPKT[1599]     = 80'hC03F7420756C74726963;
        inPKT[1600]     = 80'hC040657320706F737565;
        inPKT[1601]     = 80'hC041726520637562696C;
        inPKT[1602]     = 80'hC0426961204375726165;
        inPKT[1603]     = 80'hC0433B20437572616269;
        inPKT[1604]     = 80'hC0447475722066617563;
        inPKT[1605]     = 80'hC0456962757320646961;
        inPKT[1606]     = 80'hC0466D206C656F2C206E;
        inPKT[1607]     = 80'hC047656320657569736D;
        inPKT[1608]     = 80'hC0486F642073656D2065;
        inPKT[1609]     = 80'hC0496666696369747572;
        inPKT[1610]     = 80'hC04A2075742E20557420;
        inPKT[1611]     = 80'hC04B7665686963756C61;
        inPKT[1612]     = 80'hC04C2061756775652061;
        inPKT[1613]     = 80'hC04D63206C696265726F;
        inPKT[1614]     = 80'hC04E20696163756C6973;
        inPKT[1615]     = 80'hC04F2C206E656320656C;
        inPKT[1616]     = 80'hC050656966656E642065;
        inPKT[1617]     = 80'hC0517820706F7274612E;
        inPKT[1618]     = 80'hC052204D6F7262692068;
        inPKT[1619]     = 80'hC053656E647265726974;
        inPKT[1620]     = 80'hC0542067726176696461;
        inPKT[1621]     = 80'hC0552074696E63696475;
        inPKT[1622]     = 80'hC0566E742E2050726165;
        inPKT[1623]     = 80'hC05773656E7420646F6C;
        inPKT[1624]     = 80'hC0586F72206C61637573;
        inPKT[1625]     = 80'hC0592C2074656D707573;
        inPKT[1626]     = 80'hC05A206575206672696E;
        inPKT[1627]     = 80'hC05B67696C6C61207369;
        inPKT[1628]     = 80'hC05C7420616D65742C20;
        inPKT[1629]     = 80'hC05D656C656966656E64;
        inPKT[1630]     = 80'hC05E20696E206E756C6C;
        inPKT[1631]     = 80'hC05F612E204E756C6C61;
        inPKT[1632]     = 80'hC060206D6F6C6C697320;
        inPKT[1633]     = 80'hC06165676574206D6167;
        inPKT[1634]     = 80'hC0626E61206E65632068;
        inPKT[1635]     = 80'hC063656E647265726974;
        inPKT[1636]     = 80'hC0642E20416C69717561;
        inPKT[1637]     = 80'hC0656D20636F6E76616C;
        inPKT[1638]     = 80'hC0666C69732073656D20;
        inPKT[1639]     = 80'hC0677669746165207361;
        inPKT[1640]     = 80'hC0687069656E20646963;
        inPKT[1641]     = 80'hC06974756D2C20757420;
        inPKT[1642]     = 80'hC06A766573746962756C;
        inPKT[1643]     = 80'hC06B756D206C6F72656D;
        inPKT[1644]     = 80'hC06C206672696E67696C;
        inPKT[1645]     = 80'hC06D6C612E20446F6E65;
        inPKT[1646]     = 80'hC06E632074656C6C7573;
        inPKT[1647]     = 80'hC06F206C696265726F2C;
        inPKT[1648]     = 80'hC0702066657567696174;
        inPKT[1649]     = 80'hC0712075742066696E69;
        inPKT[1650]     = 80'hC072627573206E65632C;
        inPKT[1651]     = 80'hC07320616C697175616D;
        inPKT[1652]     = 80'hC0742073697420616D65;
        inPKT[1653]     = 80'hC07574206F7263692E20;
        inPKT[1654]     = 80'hC0764E756E6320737573;
        inPKT[1655]     = 80'hC0776369706974206E69;
        inPKT[1656]     = 80'hC078736C206574206F72;
        inPKT[1657]     = 80'hC0796E61726520766573;
        inPKT[1658]     = 80'hC07A746962756C756D2E;
        inPKT[1659]     = 80'hC07B204E756C6C616D20;
        inPKT[1660]     = 80'hC07C6C6F626F72746973;
        inPKT[1661]     = 80'hC07D2073617069656E20;
        inPKT[1662]     = 80'hC07E6A7573746F2C2073;
        inPKT[1663]     = 80'hC07F697420616D657420;
        inPKT[1664]     = 80'hC0806469676E69737369;
        inPKT[1665]     = 80'hC0816D206E756C6C6120;
        inPKT[1666]     = 80'hC082636F6E64696D656E;
        inPKT[1667]     = 80'hC08374756D20696E2E20;
        inPKT[1668]     = 80'hC084536564206D6F6C65;
        inPKT[1669]     = 80'hC0857374696520766F6C;
        inPKT[1670]     = 80'hC0867574706174206E69;
        inPKT[1671]     = 80'hC0877369206174206665;
        inPKT[1672]     = 80'hC088726D656E74756D2E;
        inPKT[1673]     = 80'hC089204E756C6C61206D;
        inPKT[1674]     = 80'hC08A6F6C657374696520;
        inPKT[1675]     = 80'hC08B6E69736920736564;
        inPKT[1676]     = 80'hC08C2074757270697320;
        inPKT[1677]     = 80'hC08D6D6F6C6573746965;
        inPKT[1678]     = 80'hC08E2C206E6F6E206961;
        inPKT[1679]     = 80'hC08F63756C6973206E75;
        inPKT[1680]     = 80'hC0906E63206661756369;
        inPKT[1681]     = 80'hC0916275732E2041656E;
        inPKT[1682]     = 80'hC09265616E20696E7465;
        inPKT[1683]     = 80'hC0937264756D20706861;
        inPKT[1684]     = 80'hC094726574726120636F;
        inPKT[1685]     = 80'hC0956E73656374657475;
        inPKT[1686]     = 80'hC096722E20457469616D;
        inPKT[1687]     = 80'hC097206578206F726369;
        inPKT[1688]     = 80'hC0982C20696163756C69;
        inPKT[1689]     = 80'hC09973206E6F6E206575;
        inPKT[1690]     = 80'hC09A69736D6F64206964;
        inPKT[1691]     = 80'hC09B2C20756C6C616D63;
        inPKT[1692]     = 80'hC09C6F72706572207363;
        inPKT[1693]     = 80'hC09D656C657269737175;
        inPKT[1694]     = 80'hC09E65206F64696F2E0D;
        inPKT[1695]     = 80'hC09F0A0D0A4E616D2075;
        inPKT[1696]     = 80'hC0A06C74726963657320;
        inPKT[1697]     = 80'hC0A1656C656966656E64;
        inPKT[1698]     = 80'hC0A2206469616D2C2065;
        inPKT[1699]     = 80'hC0A367657420736F6461;
        inPKT[1700]     = 80'hC0A46C65732073656D20;
        inPKT[1701]     = 80'hC0A56D61747469732061;
        inPKT[1702]     = 80'hC0A6632E205574207665;
        inPKT[1703]     = 80'hC0A76E656E6174697320;
        inPKT[1704]     = 80'hC0A86E69626820657520;
        inPKT[1705]     = 80'hC0A96C65637475732074;
        inPKT[1706]     = 80'hC0AA696E636964756E74;
        inPKT[1707]     = 80'hC0AB2064696374756D2E;
        inPKT[1708]     = 80'hC0AC20566976616D7573;
        inPKT[1709]     = 80'hC0AD2063757273757320;
        inPKT[1710]     = 80'hC0AE6175677565207175;
        inPKT[1711]     = 80'hC0AF6973206C6F626F72;
        inPKT[1712]     = 80'hC0B07469732065756973;
        inPKT[1713]     = 80'hC0B16D6F642E204E756E;
        inPKT[1714]     = 80'hC0B26320616C69717561;
        inPKT[1715]     = 80'hC0B36D206469616D2061;
        inPKT[1716]     = 80'hC0B47420616E74652066;
        inPKT[1717]     = 80'hC0B56163696C69736973;
        inPKT[1718]     = 80'hC0B6206D6178696D7573;
        inPKT[1719]     = 80'hC0B72E20457469616D20;
        inPKT[1720]     = 80'hC0B8736564206C6F7265;
        inPKT[1721]     = 80'hC0B96D206D6174746973;
        inPKT[1722]     = 80'hC0BA2C20636F6E76616C;
        inPKT[1723]     = 80'hC0BB6C69732075726E61;
        inPKT[1724]     = 80'hC0BC2076697461652C20;
        inPKT[1725]     = 80'hC0BD74656D7075732073;
        inPKT[1726]     = 80'hC0BE656D2E2056697661;
        inPKT[1727]     = 80'hC0BF6D75732065676573;
        inPKT[1728]     = 80'hC0C074617320766F6C75;
        inPKT[1729]     = 80'hC0C1747061742065726F;
        inPKT[1730]     = 80'hC0C27320657520756C74;
        inPKT[1731]     = 80'hC0C372696365732E2056;
        inPKT[1732]     = 80'hC0C46573746962756C75;
        inPKT[1733]     = 80'hC0C56D20756C6C616D63;
        inPKT[1734]     = 80'hC0C66F72706572206572;
        inPKT[1735]     = 80'hC0C76174206E756E632C;
        inPKT[1736]     = 80'hC0C8206E6F6E2068656E;
        inPKT[1737]     = 80'hC0C9647265726974206F;
        inPKT[1738]     = 80'hC0CA64696F2070656C6C;
        inPKT[1739]     = 80'hC0CB656E746573717565;
        inPKT[1740]     = 80'hC0CC2069642E20467573;
        inPKT[1741]     = 80'hC0CD63652075726E6120;
        inPKT[1742]     = 80'hC0CE697073756D2C206C;
        inPKT[1743]     = 80'hC0CF6163696E69612069;
        inPKT[1744]     = 80'hC0D06E20737573636970;
        inPKT[1745]     = 80'hC0D169742076656C2C20;
        inPKT[1746]     = 80'hC0D273656D7065722069;
        inPKT[1747]     = 80'hC0D36E206F64696F2E20;
        inPKT[1748]     = 80'hC0D450656C6C656E7465;
        inPKT[1749]     = 80'hC0D57371756520696420;
        inPKT[1750]     = 80'hC0D66E696268206E6973;
        inPKT[1751]     = 80'hC0D7692E20416C697175;
        inPKT[1752]     = 80'hC0D8616D20706F727461;
        inPKT[1753]     = 80'hC0D9206E69736C206574;
        inPKT[1754]     = 80'hC0DA2065782069616375;
        inPKT[1755]     = 80'hC0DB6C69732074726973;
        inPKT[1756]     = 80'hC0DC74697175652E2045;
        inPKT[1757]     = 80'hC0DD7469616D206D6173;
        inPKT[1758]     = 80'hC0DE7361206F7263692C;
        inPKT[1759]     = 80'hC0DF2065676573746173;
        inPKT[1760]     = 80'hC0E020736564206C6F72;
        inPKT[1761]     = 80'hC0E1656D20717569732C;
        inPKT[1762]     = 80'hC0E2206469676E697373;
        inPKT[1763]     = 80'hC0E3696D2073656D7065;
        inPKT[1764]     = 80'hC0E47220616E74652E20;
        inPKT[1765]     = 80'hC0E553757370656E6469;
        inPKT[1766]     = 80'hC0E67373652074696E63;
        inPKT[1767]     = 80'hC0E76964756E74206E69;
        inPKT[1768]     = 80'hC0E873692065782C2073;
        inPKT[1769]     = 80'hC0E9656420766F6C7574;
        inPKT[1770]     = 80'hC0EA7061742065737420;
        inPKT[1771]     = 80'hC0EB7661726975732076;
        inPKT[1772]     = 80'hC0EC697461652E0D0A0D;
        inPKT[1773]     = 80'hC0ED0A5365642073656D;
        inPKT[1774]     = 80'hC0EE706572206C616369;
        inPKT[1775]     = 80'hC0EF6E696120646F6C6F;
        inPKT[1776]     = 80'hC0F0722E204E616D2075;
        inPKT[1777]     = 80'hC0F1742076656C697420;
        inPKT[1778]     = 80'hC0F2696E206C61637573;
        inPKT[1779]     = 80'hC0F320636F6E73656374;
        inPKT[1780]     = 80'hC0F46574757220636F6E;
        inPKT[1781]     = 80'hC0F576616C6C69732070;
        inPKT[1782]     = 80'hC0F6656C6C656E746573;
        inPKT[1783]     = 80'hC0F77175652073656420;
        inPKT[1784]     = 80'hC0F873656D2E20537573;
        inPKT[1785]     = 80'hC0F970656E6469737365;
        inPKT[1786]     = 80'hC0FA20636F6E64696D65;
        inPKT[1787]     = 80'hC0FB6E74756D20612065;
        inPKT[1788]     = 80'hC0FC726F732069642075;
        inPKT[1789]     = 80'hC0FD6C6C616D636F7270;
        inPKT[1790]     = 80'hC0FE65722E204D6F7262;
        inPKT[1791]     = 80'hC0FF69206C7563747573;
        inPKT[1792]     = 80'hC0002075726E61207369;
        inPKT[1793]     = 80'hC0017420616D65742065;
        inPKT[1794]     = 80'hC0027569736D6F642069;
        inPKT[1795]     = 80'hC0036163756C69732E20;
        inPKT[1796]     = 80'hC00450656C6C656E7465;
        inPKT[1797]     = 80'hC0057371756520666163;
        inPKT[1798]     = 80'hC006696C69736973206D;
        inPKT[1799]     = 80'hC0076175726973206575;
        inPKT[1800]     = 80'hC00820656C656D656E74;
        inPKT[1801]     = 80'hC009756D207661726975;
        inPKT[1802]     = 80'hC00A732E204F72636920;
        inPKT[1803]     = 80'hC00B766172697573206E;
        inPKT[1804]     = 80'hC00C61746F7175652070;
        inPKT[1805]     = 80'hC00D656E617469627573;
        inPKT[1806]     = 80'hC00E206574206D61676E;
        inPKT[1807]     = 80'hC00F6973206469732070;
        inPKT[1808]     = 80'hC010617274757269656E;
        inPKT[1809]     = 80'hC01174206D6F6E746573;
        inPKT[1810]     = 80'hC0122C206E6173636574;
        inPKT[1811]     = 80'hC0137572207269646963;
        inPKT[1812]     = 80'hC014756C7573206D7573;
        inPKT[1813]     = 80'hC0152E20446F6E656320;
        inPKT[1814]     = 80'hC0166469676E69737369;
        inPKT[1815]     = 80'hC0176D20612069707375;
        inPKT[1816]     = 80'hC0186D20756C74726963;
        inPKT[1817]     = 80'hC0196965732076656E65;
        inPKT[1818]     = 80'hC01A6E617469732E2056;
        inPKT[1819]     = 80'hC01B6976616D7573206E;
        inPKT[1820]     = 80'hC01C756E632076656C69;
        inPKT[1821]     = 80'hC01D742C207665686963;
        inPKT[1822]     = 80'hC01E756C612076697461;
        inPKT[1823]     = 80'hC01F65206D6173736120;
        inPKT[1824]     = 80'hC02075742C20636F6E76;
        inPKT[1825]     = 80'hC021616C6C697320636F;
        inPKT[1826]     = 80'hC0226E73656374657475;
        inPKT[1827]     = 80'hC0237220746F72746F72;
        inPKT[1828]     = 80'hC0242E20517569737175;
        inPKT[1829]     = 80'hC0256520616C69717561;
        inPKT[1830]     = 80'hC0266D2C206E69736C20;
        inPKT[1831]     = 80'hC027636F6E6775652062;
        inPKT[1832]     = 80'hC0286C616E6469742075;
        inPKT[1833]     = 80'hC0296C74726963696573;
        inPKT[1834]     = 80'hC02A2C2075726E612074;
        inPKT[1835]     = 80'hC02B7572706973206D61;
        inPKT[1836]     = 80'hC02C74746973206D6167;
        inPKT[1837]     = 80'hC02D6E612C206E6F6E20;
        inPKT[1838]     = 80'hC02E6665726D656E7475;
        inPKT[1839]     = 80'hC02F6D20647569207665;
        inPKT[1840]     = 80'hC0306C69742065752071;
        inPKT[1841]     = 80'hC03175616D2E0D0A0D0A;
        inPKT[1842]     = 80'hC032496E207068617265;
        inPKT[1843]     = 80'hC0337472612076656C69;
        inPKT[1844]     = 80'hC0347420646F6C6F722C;
        inPKT[1845]     = 80'hC0352076697461652063;
        inPKT[1846]     = 80'hC0367572737573206F72;
        inPKT[1847]     = 80'hC03763692066696E6962;
        inPKT[1848]     = 80'hC03875732074696E6369;
        inPKT[1849]     = 80'hC03964756E742E205669;
        inPKT[1850]     = 80'hC03A76616D7573206964;
        inPKT[1851]     = 80'hC03B20746F72746F7220;
        inPKT[1852]     = 80'hC03C72686F6E6375732C;
        inPKT[1853]     = 80'hC03D2073616769747469;
        inPKT[1854]     = 80'hC03E73206469616D2065;
        inPKT[1855]     = 80'hC03F6765742C20707265;
        inPKT[1856]     = 80'hC0407469756D206D6175;
        inPKT[1857]     = 80'hC0417269732E20506861;
        inPKT[1858]     = 80'hC04273656C6C75732065;
        inPKT[1859]     = 80'hC0436C656D656E74756D;
        inPKT[1860]     = 80'hC04420656E696D206665;
        inPKT[1861]     = 80'hC0456C69732E204D6175;
        inPKT[1862]     = 80'hC046726973206575206E;
        inPKT[1863]     = 80'hC0476571756520656765;
        inPKT[1864]     = 80'hC0487420707572757320;
        inPKT[1865]     = 80'hC04968656E6472657269;
        inPKT[1866]     = 80'hC04A7420677261766964;
        inPKT[1867]     = 80'hC04B612E20416C697175;
        inPKT[1868]     = 80'hC04C616D206C69626572;
        inPKT[1869]     = 80'hC04D6F206E6962682C20;
        inPKT[1870]     = 80'hC04E636F6E76616C6C69;
        inPKT[1871]     = 80'hC04F732061206E69736C;
        inPKT[1872]     = 80'hC0502065742C2068656E;
        inPKT[1873]     = 80'hC0516472657269742076;
        inPKT[1874]     = 80'hC0526573746962756C75;
        inPKT[1875]     = 80'hC0536D2066656C69732E;
        inPKT[1876]     = 80'hC05420446F6E65632065;
        inPKT[1877]     = 80'hC0557569736D6F642066;
        inPKT[1878]     = 80'hC05665726D656E74756D;
        inPKT[1879]     = 80'hC0572074757270697320;
        inPKT[1880]     = 80'hC058657520617563746F;
        inPKT[1881]     = 80'hC059722E2041656E6561;
        inPKT[1882]     = 80'hC05A6E20626962656E64;
        inPKT[1883]     = 80'hC05B756D207475727069;
        inPKT[1884]     = 80'hC05C7320696E206F6469;
        inPKT[1885]     = 80'hC05D6F20636F6E76616C;
        inPKT[1886]     = 80'hC05E6C69732C20766974;
        inPKT[1887]     = 80'hC05F6165207661726975;
        inPKT[1888]     = 80'hC06073206578206C616F;
        inPKT[1889]     = 80'hC061726565742E204675;
        inPKT[1890]     = 80'hC0627363652076656C20;
        inPKT[1891]     = 80'hC0636D69207669746165;
        inPKT[1892]     = 80'hC06420646F6C6F722066;
        inPKT[1893]     = 80'hC0656575676961742076;
        inPKT[1894]     = 80'hC066756C707574617465;
        inPKT[1895]     = 80'hC067206E656320757420;
        inPKT[1896]     = 80'hC0686E756E632E204372;
        inPKT[1897]     = 80'hC0696173206461706962;
        inPKT[1898]     = 80'hC06A75732C20616E7465;
        inPKT[1899]     = 80'hC06B2069642076656869;
        inPKT[1900]     = 80'hC06C63756C6120616C69;
        inPKT[1901]     = 80'hC06D7175616D2C20656C;
        inPKT[1902]     = 80'hC06E69742065726F7320;
        inPKT[1903]     = 80'hC06F7361676974746973;
        inPKT[1904]     = 80'hC070206D692C206E6F6E;
        inPKT[1905]     = 80'hC07120656C656966656E;
        inPKT[1906]     = 80'hC07264206578206E756C;
        inPKT[1907]     = 80'hC0736C61206567657420;
        inPKT[1908]     = 80'hC07476656C69742E2053;
        inPKT[1909]     = 80'hC075757370656E646973;
        inPKT[1910]     = 80'hC0767365206964206469;
        inPKT[1911]     = 80'hC077616D206475692E20;
        inPKT[1912]     = 80'hC07853757370656E6469;
        inPKT[1913]     = 80'hC0797373652070726574;
        inPKT[1914]     = 80'hC07A69756D206A757374;
        inPKT[1915]     = 80'hC07B6F20736564206E69;
        inPKT[1916]     = 80'hC07C626820706F727474;
        inPKT[1917]     = 80'hC07D69746F722C207665;
        inPKT[1918]     = 80'hC07E6C20696E74657264;
        inPKT[1919]     = 80'hC07F756D206D61757269;
        inPKT[1920]     = 80'hC08073206D6178696D75;
        inPKT[1921]     = 80'hC081732E20557420616C;
        inPKT[1922]     = 80'hC082697175616D206C61;
        inPKT[1923]     = 80'hC0836375732070757275;
        inPKT[1924]     = 80'hC084732C207369742061;
        inPKT[1925]     = 80'hC0856D657420696D7065;
        inPKT[1926]     = 80'hC0867264696574206E69;
        inPKT[1927]     = 80'hC0876268206665756769;
        inPKT[1928]     = 80'hC08861742069642E2049;
        inPKT[1929]     = 80'hC0896E7465676572206C;
        inPKT[1930]     = 80'hC08A6F72656D206D6175;
        inPKT[1931]     = 80'hC08B7269732C20707265;
        inPKT[1932]     = 80'hC08C7469756D206E6F6E;
        inPKT[1933]     = 80'hC08D206E697369206574;
        inPKT[1934]     = 80'hC08E2C20646170696275;
        inPKT[1935]     = 80'hC08F732066696E696275;
        inPKT[1936]     = 80'hC09073206F7263692E0D;
        inPKT[1937]     = 80'hC0910A0D0A5665737469;
        inPKT[1938]     = 80'hC09262756C756D206961;
        inPKT[1939]     = 80'hC09363756C69732C206D;
        inPKT[1940]     = 80'hC09461676E6120617420;
        inPKT[1941]     = 80'hC0956D6174746973206D;
        inPKT[1942]     = 80'hC0966178696D75732C20;
        inPKT[1943]     = 80'hC0976172637520657261;
        inPKT[1944]     = 80'hC0987420646170696275;
        inPKT[1945]     = 80'hC09973206E756E632C20;
        inPKT[1946]     = 80'hC09A6120766172697573;
        inPKT[1947]     = 80'hC09B206D657475732066;
        inPKT[1948]     = 80'hC09C656C697320736564;
        inPKT[1949]     = 80'hC09D206F7263692E204E;
        inPKT[1950]     = 80'hC09E756C6C616D206D69;
        inPKT[1951]     = 80'hC09F206E6962682C2065;
        inPKT[1952]     = 80'hC0A06C656966656E6420;
        inPKT[1953]     = 80'hC0A16E656320756C7472;
        inPKT[1954]     = 80'hC0A269636573206E6563;
        inPKT[1955]     = 80'hC0A32C20636F6E736563;
        inPKT[1956]     = 80'hC0A47465747572206163;
        inPKT[1957]     = 80'hC0A520656E696D2E2053;
        inPKT[1958]     = 80'hC0A66564206C75637475;
        inPKT[1959]     = 80'hC0A7732073656D207175;
        inPKT[1960]     = 80'hC0A869732074656D706F;
        inPKT[1961]     = 80'hC0A97220636F6E677565;
        inPKT[1962]     = 80'hC0AA2E2053757370656E;
        inPKT[1963]     = 80'hC0AB646973736520706F;
        inPKT[1964]     = 80'hC0AC74656E74692E2045;
        inPKT[1965]     = 80'hC0AD7469616D20656765;
        inPKT[1966]     = 80'hC0AE74206C696265726F;
        inPKT[1967]     = 80'hC0AF2076656C69742E20;
        inPKT[1968]     = 80'hC0B04475697320766573;
        inPKT[1969]     = 80'hC0B1746962756C756D20;
        inPKT[1970]     = 80'hC0B2636F6E7365717561;
        inPKT[1971]     = 80'hC0B37420706F7274612E;
        inPKT[1972]     = 80'hC0B4204D617572697320;
        inPKT[1973]     = 80'hC0B5706F72747469746F;
        inPKT[1974]     = 80'hC0B67220747572706973;
        inPKT[1975]     = 80'hC0B720696E206D617373;
        inPKT[1976]     = 80'hC0B86120616C69717561;
        inPKT[1977]     = 80'hC0B96D20636F6E677565;
        inPKT[1978]     = 80'hC0BA2E204E756C6C6120;
        inPKT[1979]     = 80'hC0BB636F6E7365637465;
        inPKT[1980]     = 80'hC0BC7475722075726E61;
        inPKT[1981]     = 80'hC0BD206D657475732C20;
        inPKT[1982]     = 80'hC0BE696420696163756C;
        inPKT[1983]     = 80'hC0BF6973206E756E6320;
        inPKT[1984]     = 80'hC0C0756C747269636965;
        inPKT[1985]     = 80'hC0C17320656765742E20;
        inPKT[1986]     = 80'hC0C24375726162697475;
        inPKT[1987]     = 80'hC0C372206D6175726973;
        inPKT[1988]     = 80'hC0C4206E657175652C20;
        inPKT[1989]     = 80'hC0C5626962656E64756D;
        inPKT[1990]     = 80'hC0C6207365642065726F;
        inPKT[1991]     = 80'hC0C7732061742C206D61;
        inPKT[1992]     = 80'hC0C878696D757320756C;
        inPKT[1993]     = 80'hC0C97472696365732074;
        inPKT[1994]     = 80'hC0CA75727069732E0D0A;
        inPKT[1995]     = 80'hC0CB496E74657264756D;
        inPKT[1996]     = 80'hC0CC206574206D616C65;
        inPKT[1997]     = 80'hC0CD7375616461206661;
        inPKT[1998]     = 80'hC0CE6D65732061632061;
        inPKT[1999]     = 80'hC0CF6E74652069707375;
        inPKT[2000]     = 80'hC0D06D207072696D6973;
        inPKT[2001]     = 80'hC0D120696E2066617563;
        inPKT[2002]     = 80'hC0D2696275732E205065;
        inPKT[2003]     = 80'hC0D36C6C656E74657371;
        inPKT[2004]     = 80'hC0D4756520736F6C6C69;
        inPKT[2005]     = 80'hC0D56369747564696E20;
        inPKT[2006]     = 80'hC0D6626C616E64697420;
        inPKT[2007]     = 80'hC0D76665726D656E7475;
        inPKT[2008]     = 80'hC0D86D2E2050656C6C65;
        inPKT[2009]     = 80'hC0D96E74657371756520;
        inPKT[2010]     = 80'hC0DA6E6F6E206C696775;
        inPKT[2011]     = 80'hC0DB6C61206575206572;
        inPKT[2012]     = 80'hC0DC61742076656E656E;
        inPKT[2013]     = 80'hC0DD6174697320657569;
        inPKT[2014]     = 80'hC0DE736D6F642E205065;
        inPKT[2015]     = 80'hC0DF6C6C656E74657371;
        inPKT[2016]     = 80'hC0E0756520736F64616C;
        inPKT[2017]     = 80'hC0E16573207665737469;
        inPKT[2018]     = 80'hC0E262756C756D20636F;
        inPKT[2019]     = 80'hC0E36E76616C6C69732E;
        inPKT[2020]     = 80'hC0E42050726F696E206D;
        inPKT[2021]     = 80'hC0E56F6C657374696520;
        inPKT[2022]     = 80'hC0E67072657469756D20;
        inPKT[2023]     = 80'hC0E765726F732076656C;
        inPKT[2024]     = 80'hC0E82065676573746173;
        inPKT[2025]     = 80'hC0E92E204D6F72626920;
        inPKT[2026]     = 80'hC0EA736F6C6C69636974;
        inPKT[2027]     = 80'hC0EB7564696E20707572;
        inPKT[2028]     = 80'hC0EC7573206163206665;
        inPKT[2029]     = 80'hC0ED726D656E74756D20;
        inPKT[2030]     = 80'hC0EE6D61747469732E20;
        inPKT[2031]     = 80'hC0EF4E756E632076656C;
        inPKT[2032]     = 80'hC0F02074696E63696475;
        inPKT[2033]     = 80'hC0F16E74206C69626572;
        inPKT[2034]     = 80'hC0F26F2E204E756C6C61;
        inPKT[2035]     = 80'hC0F320616C6971756574;
        inPKT[2036]     = 80'hC0F420697073756D206E;
        inPKT[2037]     = 80'hC0F56563207175616D20;
        inPKT[2038]     = 80'hC0F6696D706572646965;
        inPKT[2039]     = 80'hC0F77420696E74657264;
        inPKT[2040]     = 80'hC0F8756D2E2050726165;
        inPKT[2041]     = 80'hC0F973656E74206C6967;
        inPKT[2042]     = 80'hC0FA756C612066656C69;
        inPKT[2043]     = 80'hC0FB732C20696163756C;
        inPKT[2044]     = 80'hC0FC697320617420616C;
        inPKT[2045]     = 80'hC0FD6971756574206174;
        inPKT[2046]     = 80'hC0FE2C20736167697474;
        inPKT[2047]     = 80'hC0FF6973207175697320;
        inPKT[2048]     = 80'hC000656C69742E0D0A51;
        inPKT[2049]     = 80'hC0017569737175652076;
        inPKT[2050]     = 80'hC002656C20696D706572;
        inPKT[2051]     = 80'hC00364696574206E6962;
        inPKT[2052]     = 80'hC004682E205068617365;
        inPKT[2053]     = 80'hC0056C6C757320727574;
        inPKT[2054]     = 80'hC00672756D206469676E;
        inPKT[2055]     = 80'hC007697373696D207269;
        inPKT[2056]     = 80'hC008737573206E6F6E20;
        inPKT[2057]     = 80'hC00974696E636964756E;
        inPKT[2058]     = 80'hC00A742E205665737469;
        inPKT[2059]     = 80'hC00B62756C756D206E75;
        inPKT[2060]     = 80'hC00C6E6320697073756D;
        inPKT[2061]     = 80'hC00D2C2076656E656E61;
        inPKT[2062]     = 80'hC00E7469732065676574;
        inPKT[2063]     = 80'hC00F20706F7274612069;
        inPKT[2064]     = 80'hC0106E2C20636F6E7365;
        inPKT[2065]     = 80'hC0116374657475722065;
        inPKT[2066]     = 80'hC0127520657261742E20;
        inPKT[2067]     = 80'hC013446F6E6563207665;
        inPKT[2068]     = 80'hC014686963756C612061;
        inPKT[2069]     = 80'hC0156E74652076656C20;
        inPKT[2070]     = 80'hC01672686F6E63757320;
        inPKT[2071]     = 80'hC0176661756369627573;
        inPKT[2072]     = 80'hC0182E2050656C6C656E;
        inPKT[2073]     = 80'hC019746573717565206A;
        inPKT[2074]     = 80'hC01A7573746F20746F72;
        inPKT[2075]     = 80'hC01B746F722C20766F6C;
        inPKT[2076]     = 80'hC01C757470617420696E;
        inPKT[2077]     = 80'hC01D206D617572697320;
        inPKT[2078]     = 80'hC01E61742C2076617269;
        inPKT[2079]     = 80'hC01F7573207068617265;
        inPKT[2080]     = 80'hC0207472612072697375;
        inPKT[2081]     = 80'hC021732E205175697371;
        inPKT[2082]     = 80'hC0227565207574206469;
        inPKT[2083]     = 80'hC023616D207375736369;
        inPKT[2084]     = 80'hC0247069742C20736F6C;
        inPKT[2085]     = 80'hC0256C69636974756469;
        inPKT[2086]     = 80'hC0266E2073617069656E;
        inPKT[2087]     = 80'hC0272065742C20696E74;
        inPKT[2088]     = 80'hC028657264756D206C61;
        inPKT[2089]     = 80'hC0296375732E204D6F72;
        inPKT[2090]     = 80'hC02A6269207269737573;
        inPKT[2091]     = 80'hC02B2073656D2C207065;
        inPKT[2092]     = 80'hC02C6C6C656E74657371;
        inPKT[2093]     = 80'hC02D7565206574207475;
        inPKT[2094]     = 80'hC02E7270697320696E2C;
        inPKT[2095]     = 80'hC02F20626C616E646974;
        inPKT[2096]     = 80'hC03020736F6C6C696369;
        inPKT[2097]     = 80'hC031747564696E207365;
        inPKT[2098]     = 80'hC0326D2E205365642065;
        inPKT[2099]     = 80'hC0336666696369747572;
        inPKT[2100]     = 80'hC034206C696265726F20;
        inPKT[2101]     = 80'hC0357175697320707265;
        inPKT[2102]     = 80'hC0367469756D20707265;
        inPKT[2103]     = 80'hC0377469756D2E204E75;
        inPKT[2104]     = 80'hC0386C6C616D20617563;
        inPKT[2105]     = 80'hC039746F722073616769;
        inPKT[2106]     = 80'hC03A74746973206C6F72;
        inPKT[2107]     = 80'hC03B656D2C2061632075;
        inPKT[2108]     = 80'hC03C6C74726963657320;
        inPKT[2109]     = 80'hC03D61726375206D6178;
        inPKT[2110]     = 80'hC03E696D757320656765;
        inPKT[2111]     = 80'hC03F742E0D0A56657374;
        inPKT[2112]     = 80'hC0406962756C756D2076;
        inPKT[2113]     = 80'hC0416F6C757470617420;
        inPKT[2114]     = 80'hC0426C6967756C612061;
        inPKT[2115]     = 80'hC0437563746F72207365;
        inPKT[2116]     = 80'hC0446D20766976657272;
        inPKT[2117]     = 80'hC045612C20756C6C616D;
        inPKT[2118]     = 80'hC046636F727065722065;
        inPKT[2119]     = 80'hC0477569736D6F64206E;
        inPKT[2120]     = 80'hC0486571756520706F72;
        inPKT[2121]     = 80'hC049747469746F722E20;
        inPKT[2122]     = 80'hC04A53757370656E6469;
        inPKT[2123]     = 80'hC04B7373652076697665;
        inPKT[2124]     = 80'hC04C727261207363656C;
        inPKT[2125]     = 80'hC04D6572697371756520;
        inPKT[2126]     = 80'hC04E6F64696F2072686F;
        inPKT[2127]     = 80'hC04F6E63757320766F6C;
        inPKT[2128]     = 80'hC05075747061742E2041;
        inPKT[2129]     = 80'hC0516C697175616D2065;
        inPKT[2130]     = 80'hC05272617420766F6C75;
        inPKT[2131]     = 80'hC053747061742E205375;
        inPKT[2132]     = 80'hC0547370656E64697373;
        inPKT[2133]     = 80'hC0556520706F74656E74;
        inPKT[2134]     = 80'hC056692E20496E206861;
        inPKT[2135]     = 80'hC0576320686162697461;
        inPKT[2136]     = 80'hC05873736520706C6174;
        inPKT[2137]     = 80'hC0596561206469637475;
        inPKT[2138]     = 80'hC05A6D73742E2050726F;
        inPKT[2139]     = 80'hC05B696E207574206E75;
        inPKT[2140]     = 80'hC05C6C6C612075742064;
        inPKT[2141]     = 80'hC05D7569207363656C65;
        inPKT[2142]     = 80'hC05E7269737175652064;
        inPKT[2143]     = 80'hC05F696374756D2E2051;
        inPKT[2144]     = 80'hC0607569737175652073;
        inPKT[2145]     = 80'hC0617573636970697420;
        inPKT[2146]     = 80'hC0626E69626820706F73;
        inPKT[2147]     = 80'hC0637565726520717561;
        inPKT[2148]     = 80'hC0646D2076756C707574;
        inPKT[2149]     = 80'hC0656174652C20657520;
        inPKT[2150]     = 80'hC0666C6163696E696120;
        inPKT[2151]     = 80'hC067616E746520677261;
        inPKT[2152]     = 80'hC068766964612E204375;
        inPKT[2153]     = 80'hC0697261626974757220;
        inPKT[2154]     = 80'hC06A6D61737361206C6F;
        inPKT[2155]     = 80'hC06B72656D2C206F726E;
        inPKT[2156]     = 80'hC06C617265206575206D;
        inPKT[2157]     = 80'hC06D6F6C6C6973206174;
        inPKT[2158]     = 80'hC06E2C20706861726574;
        inPKT[2159]     = 80'hC06F7261206E6563206D;
        inPKT[2160]     = 80'hC070617373612E204E75;
        inPKT[2161]     = 80'hC0716C6C612066696E69;
        inPKT[2162]     = 80'hC07262757320656C6569;
        inPKT[2163]     = 80'hC07366656E64206F7263;
        inPKT[2164]     = 80'hC074692073697420616D;
        inPKT[2165]     = 80'hC075657420636F6E7365;
        inPKT[2166]     = 80'hC0766374657475722E20;
        inPKT[2167]     = 80'hC0775365642074656D70;
        inPKT[2168]     = 80'hC0787573207669746165;
        inPKT[2169]     = 80'hC0792061726375206E65;
        inPKT[2170]     = 80'hC07A63206665726D656E;
        inPKT[2171]     = 80'hC07B74756D2E2041656E;
        inPKT[2172]     = 80'hC07C65616E2070656C6C;
        inPKT[2173]     = 80'hC07D656E746573717565;
        inPKT[2174]     = 80'hC07E2076697461652064;
        inPKT[2175]     = 80'hC07F6F6C6F7220696E20;
        inPKT[2176]     = 80'hC080616363756D73616E;
        inPKT[2177]     = 80'hC0812E20437261732064;
        inPKT[2178]     = 80'hC08269676E697373696D;
        inPKT[2179]     = 80'hC0832076756C70757461;
        inPKT[2180]     = 80'hC0847465206D6F6C6C69;
        inPKT[2181]     = 80'hC085732E204D61757269;
        inPKT[2182]     = 80'hC0867320706F72746120;
        inPKT[2183]     = 80'hC08776656E656E617469;
        inPKT[2184]     = 80'hC088732072697375732C;
        inPKT[2185]     = 80'hC0892065752074726973;
        inPKT[2186]     = 80'hC08A746971756520646F;
        inPKT[2187]     = 80'hC08B6C6F722072757472;
        inPKT[2188]     = 80'hC08C756D20696E2E2046;
        inPKT[2189]     = 80'hC08D7573636520636F6E;
        inPKT[2190]     = 80'hC08E64696D656E74756D;
        inPKT[2191]     = 80'hC08F206F726369206665;
        inPKT[2192]     = 80'hC0906C69732C20736974;
        inPKT[2193]     = 80'hC09120616D657420636F;
        inPKT[2194]     = 80'hC0926E76616C6C697320;
        inPKT[2195]     = 80'hC0936C696265726F2074;
        inPKT[2196]     = 80'hC094696E636964756E74;
        inPKT[2197]     = 80'hC0952061632E0D0A5665;
        inPKT[2198]     = 80'hC09673746962756C756D;
        inPKT[2199]     = 80'hC09720696D7065726469;
        inPKT[2200]     = 80'hC098657420656C697420;
        inPKT[2201]     = 80'hC09974656D706F722071;
        inPKT[2202]     = 80'hC09A75616D2067726176;
        inPKT[2203]     = 80'hC09B6964612C20757420;
        inPKT[2204]     = 80'hC09C6D616C6573756164;
        inPKT[2205]     = 80'hC09D612074656C6C7573;
        inPKT[2206]     = 80'hC09E20696D7065726469;
        inPKT[2207]     = 80'hC09F65742E2050686173;
        inPKT[2208]     = 80'hC0A0656C6C7573206F64;
        inPKT[2209]     = 80'hC0A1696F2073656D2C20;
        inPKT[2210]     = 80'hC0A26D61747469732073;
        inPKT[2211]     = 80'hC0A3656420756C747269;
        inPKT[2212]     = 80'hC0A46365732061742C20;
        inPKT[2213]     = 80'hC0A57669766572726120;
        inPKT[2214]     = 80'hC0A676656C206475692E;
        inPKT[2215]     = 80'hC0A7204E756E63207572;
        inPKT[2216]     = 80'hC0A86E61206D65747573;
        inPKT[2217]     = 80'hC0A92C206C7563747573;
        inPKT[2218]     = 80'hC0AA206163206D617869;
        inPKT[2219]     = 80'hC0AB6D757320696E2C20;
        inPKT[2220]     = 80'hC0AC636F6E7365637465;
        inPKT[2221]     = 80'hC0AD747572206E6F6E20;
        inPKT[2222]     = 80'hC0AE6E6973692E204E75;
        inPKT[2223]     = 80'hC0AF6C6C612073697420;
        inPKT[2224]     = 80'hC0B0616D657420626962;
        inPKT[2225]     = 80'hC0B1656E64756D207665;
        inPKT[2226]     = 80'hC0B26C69742E20446F6E;
        inPKT[2227]     = 80'hC0B36563207175697320;
        inPKT[2228]     = 80'hC0B4656E696D206E6F6E;
        inPKT[2229]     = 80'hC0B52072697375732062;
        inPKT[2230]     = 80'hC0B66C616E6469742066;
        inPKT[2231]     = 80'hC0B76163696C69736973;
        inPKT[2232]     = 80'hC0B82071756973206E65;
        inPKT[2233]     = 80'hC0B9632072697375732E;
        inPKT[2234]     = 80'hC0BA2043757261626974;
        inPKT[2235]     = 80'hC0BB7572206575206573;
        inPKT[2236]     = 80'hC0BC7420766974616520;
        inPKT[2237]     = 80'hC0BD6C65637475732062;
        inPKT[2238]     = 80'hC0BE6C616E6469742061;
        inPKT[2239]     = 80'hC0BF6C69717565742E20;
        inPKT[2240]     = 80'hC0C0566573746962756C;
        inPKT[2241]     = 80'hC0C1756D20616E746520;
        inPKT[2242]     = 80'hC0C2697073756D207072;
        inPKT[2243]     = 80'hC0C3696D697320696E20;
        inPKT[2244]     = 80'hC0C46661756369627573;
        inPKT[2245]     = 80'hC0C5206F726369206C75;
        inPKT[2246]     = 80'hC0C66374757320657420;
        inPKT[2247]     = 80'hC0C7756C747269636573;
        inPKT[2248]     = 80'hC0C820706F7375657265;
        inPKT[2249]     = 80'hC0C920637562696C6961;
        inPKT[2250]     = 80'hC0CA2043757261653B20;
        inPKT[2251]     = 80'hC0CB566573746962756C;
        inPKT[2252]     = 80'hC0CC756D206163206469;
        inPKT[2253]     = 80'hC0CD676E697373696D20;
        inPKT[2254]     = 80'hC0CE6E756E632E205175;
        inPKT[2255]     = 80'hC0CF697371756520696E;
        inPKT[2256]     = 80'hC0D02073616769747469;
        inPKT[2257]     = 80'hC0D1732074656C6C7573;
        inPKT[2258]     = 80'hC0D22C2073697420616D;
        inPKT[2259]     = 80'hC0D36574206665726D65;
        inPKT[2260]     = 80'hC0D46E74756D206E6962;
        inPKT[2261]     = 80'hC0D5682E0D0A496E2064;
        inPKT[2262]     = 80'hC0D669676E697373696D;
        inPKT[2263]     = 80'hC0D72072697375732076;
        inPKT[2264]     = 80'hC0D86974616520707572;
        inPKT[2265]     = 80'hC0D97573207665737469;
        inPKT[2266]     = 80'hC0DA62756C756D2C2061;
        inPKT[2267]     = 80'hC0DB7420656C656D656E;
        inPKT[2268]     = 80'hC0DC74756D206E756C6C;
        inPKT[2269]     = 80'hC0DD6120706F73756572;
        inPKT[2270]     = 80'hC0DE652E20536564206D;
        inPKT[2271]     = 80'hC0DF6174746973206E75;
        inPKT[2272]     = 80'hC0E06E63206E6962682E;
        inPKT[2273]     = 80'hC0E12053757370656E64;
        inPKT[2274]     = 80'hC0E2697373652070656C;
        inPKT[2275]     = 80'hC0E36C656E7465737175;
        inPKT[2276]     = 80'hC0E46520706C61636572;
        inPKT[2277]     = 80'hC0E56174207363656C65;
        inPKT[2278]     = 80'hC0E67269737175652E20;
        inPKT[2279]     = 80'hC0E741656E65616E2066;
        inPKT[2280]     = 80'hC0E8657567696174206D;
        inPKT[2281]     = 80'hC0E96175726973206964;
        inPKT[2282]     = 80'hC0EA20636F6E67756520;
        inPKT[2283]     = 80'hC0EB6C6163696E69612E;
        inPKT[2284]     = 80'hC0EC20457469616D2073;
        inPKT[2285]     = 80'hC0ED7573636970697420;
        inPKT[2286]     = 80'hC0EE6C6967756C612074;
        inPKT[2287]     = 80'hC0EF656C6C75732C2061;
        inPKT[2288]     = 80'hC0F020636F6E67756520;
        inPKT[2289]     = 80'hC0F16C65637475732061;
        inPKT[2290]     = 80'hC0F26C697175616D2076;
        inPKT[2291]     = 80'hC0F365686963756C612E;
        inPKT[2292]     = 80'hC0F42053757370656E64;
        inPKT[2293]     = 80'hC0F56973736520656765;
        inPKT[2294]     = 80'hC0F67420616E74652076;
        inPKT[2295]     = 80'hC0F7656C20656E696D20;
        inPKT[2296]     = 80'hC0F86D616C6573756164;
        inPKT[2297]     = 80'hC0F96120766976657272;
        inPKT[2298]     = 80'hC0FA612E2050726F696E;
        inPKT[2299]     = 80'hC0FB2074696E63696475;
        inPKT[2300]     = 80'hC0FC6E74206172637520;
        inPKT[2301]     = 80'hC0FD656765742076756C;
        inPKT[2302]     = 80'hC0FE7075746174652061;
        inPKT[2303]     = 80'hC0FF6363756D73616E2E;
        inPKT[2304]     = 80'hC00020496E2076697461;
        inPKT[2305]     = 80'hC00165206469616D206E;
        inPKT[2306]     = 80'hC0026962682E204D6F72;
        inPKT[2307]     = 80'hC0036269206D6178696D;
        inPKT[2308]     = 80'hC00475732066656C6973;
        inPKT[2309]     = 80'hC00520696420636F6E73;
        inPKT[2310]     = 80'hC0066563746574757220;
        inPKT[2311]     = 80'hC007616C697175616D2E;
        inPKT[2312]     = 80'hC008204E756C6C612066;
        inPKT[2313]     = 80'hC0096163696C6973692E;
        inPKT[2314]     = 80'hC00A0D0A566573746962;
        inPKT[2315]     = 80'hC00B756C756D20766573;
        inPKT[2316]     = 80'hC00C746962756C756D20;
        inPKT[2317]     = 80'hC00D6566666963697475;
        inPKT[2318]     = 80'hC00E7220746F72746F72;
        inPKT[2319]     = 80'hC00F2073697420616D65;
        inPKT[2320]     = 80'hC0107420666163696C69;
        inPKT[2321]     = 80'hC0117369732E204D6165;
        inPKT[2322]     = 80'hC01263656E6173206E6F;
        inPKT[2323]     = 80'hC0136E2074656C6C7573;
        inPKT[2324]     = 80'hC014206F7263692E2050;
        inPKT[2325]     = 80'hC015686173656C6C7573;
        inPKT[2326]     = 80'hC016206E6F6E206C7563;
        inPKT[2327]     = 80'hC017747573206A757374;
        inPKT[2328]     = 80'hC0186F2C206174207375;
        inPKT[2329]     = 80'hC0197363697069742074;
        inPKT[2330]     = 80'hC01A656C6C75732E2046;
        inPKT[2331]     = 80'hC01B757363652068656E;
        inPKT[2332]     = 80'hC01C647265726974206E;
        inPKT[2333]     = 80'hC01D6563206E69626820;
        inPKT[2334]     = 80'hC01E76656C2063757273;
        inPKT[2335]     = 80'hC01F75732E2053757370;
        inPKT[2336]     = 80'hC020656E646973736520;
        inPKT[2337]     = 80'hC021706F74656E74692E;
        inPKT[2338]     = 80'hC0222044756973206C69;
        inPKT[2339]     = 80'hC02367756C612066656C;
        inPKT[2340]     = 80'hC02469732C2065666669;
        inPKT[2341]     = 80'hC0256369747572206574;
        inPKT[2342]     = 80'hC0262076656C69742061;
        inPKT[2343]     = 80'hC027742C20666163696C;
        inPKT[2344]     = 80'hC0286973697320636F6E;
        inPKT[2345]     = 80'hC02976616C6C6973206A;
        inPKT[2346]     = 80'hC02A7573746F2E204E75;
        inPKT[2347]     = 80'hC02B6C6C616D206C6F62;
        inPKT[2348]     = 80'hC02C6F72746973207065;
        inPKT[2349]     = 80'hC02D6C6C656E74657371;
        inPKT[2350]     = 80'hC02E756520736F6C6C69;
        inPKT[2351]     = 80'hC02F6369747564696E2E;
        inPKT[2352]     = 80'hC030204E616D20736974;
        inPKT[2353]     = 80'hC03120616D657420646F;
        inPKT[2354]     = 80'hC0326C6F722073697420;
        inPKT[2355]     = 80'hC033616D6574206C6563;
        inPKT[2356]     = 80'hC03474757320696D7065;
        inPKT[2357]     = 80'hC035726469657420636F;
        inPKT[2358]     = 80'hC0366E7365717561742E;
        inPKT[2359]     = 80'hC03720416C697175616D;
        inPKT[2360]     = 80'hC038206C756374757320;
        inPKT[2361]     = 80'hC0397363656C65726973;
        inPKT[2362]     = 80'hC03A7175652070757275;
        inPKT[2363]     = 80'hC03B732C206964206672;
        inPKT[2364]     = 80'hC03C696E67696C6C6120;
        inPKT[2365]     = 80'hC03D73656D20766F6C75;
        inPKT[2366]     = 80'hC03E747061742061632E;
        inPKT[2367]     = 80'hC03F205365642074656D;
        inPKT[2368]     = 80'hC040706F722C20656E69;
        inPKT[2369]     = 80'hC0416D20656765742065;
        inPKT[2370]     = 80'hC0427569736D6F642066;
        inPKT[2371]     = 80'hC0436163696C69736973;
        inPKT[2372]     = 80'hC0442C206E6973692065;
        inPKT[2373]     = 80'hC045782073656D706572;
        inPKT[2374]     = 80'hC04620697073756D2C20;
        inPKT[2375]     = 80'hC047696E207361676974;
        inPKT[2376]     = 80'hC048746973206F726369;
        inPKT[2377]     = 80'hC049207175616D20696E;
        inPKT[2378]     = 80'hC04A206C65637475732E;
        inPKT[2379]     = 80'hC04B2055742076697461;
        inPKT[2380]     = 80'hC04C6520656C6974206C;
        inPKT[2381]     = 80'hC04D6967756C612E204E;
        inPKT[2382]     = 80'hC04E756E632065676573;
        inPKT[2383]     = 80'hC04F7461732C206D6920;
        inPKT[2384]     = 80'hC0507669746165206961;
        inPKT[2385]     = 80'hC05163756C6973206D61;
        inPKT[2386]     = 80'hC052747469732C206475;
        inPKT[2387]     = 80'hC05369206E6962682065;
        inPKT[2388]     = 80'hC0546C656966656E6420;
        inPKT[2389]     = 80'hC0556E69736C2C206567;
        inPKT[2390]     = 80'hC056657420706F727461;
        inPKT[2391]     = 80'hC057206C696265726F20;
        inPKT[2392]     = 80'hC0586175677565207175;
        inPKT[2393]     = 80'hC059697320656E696D2E;
        inPKT[2394]     = 80'hC05A2053656420736974;
        inPKT[2395]     = 80'hC05B20616D6574207075;
        inPKT[2396]     = 80'hC05C6C76696E61722065;
        inPKT[2397]     = 80'hC05D782C2076656C2070;
        inPKT[2398]     = 80'hC05E656C6C656E746573;
        inPKT[2399]     = 80'hC05F717565206C616375;
        inPKT[2400]     = 80'hC06073206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
