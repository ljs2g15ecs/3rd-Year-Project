`include "SIMON_defintions.svh"
