`include "SIMON_defintions.svh"

module test_SIMON_4872_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 1600
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 112'hE1001211100A0908020100000000;
        inPKT[1]        = 112'hC1014C6F72656D20697073756D20;
        inPKT[2]        = 112'hC102646F6C6F722073697420616D;
        inPKT[3]        = 112'hC10365742C20636F6E7365637465;
        inPKT[4]        = 112'hC104747572206164697069736369;
        inPKT[5]        = 112'hC1056E6720656C69742E20437572;
        inPKT[6]        = 112'hC10661626974757220756C6C616D;
        inPKT[7]        = 112'hC107636F727065722074656D7075;
        inPKT[8]        = 112'hC10873206E6973692C2065742070;
        inPKT[9]        = 112'hC1096F73756572652075726E612E;
        inPKT[10]       = 112'hC10A2041656E65616E2073656420;
        inPKT[11]       = 112'hC10B67726176696461206C616375;
        inPKT[12]       = 112'hC10C732E204E756C6C6120666163;
        inPKT[13]       = 112'hC10D696C6973692E204E756C6C61;
        inPKT[14]       = 112'hC10E2074656D707573206F726369;
        inPKT[15]       = 112'hC10F207175697320656C69742066;
        inPKT[16]       = 112'hC1106575676961742C2076656C20;
        inPKT[17]       = 112'hC11173656D706572206C656F2069;
        inPKT[18]       = 112'hC1126D706572646965742E204D61;
        inPKT[19]       = 112'hC1136563656E6173206574206E75;
        inPKT[20]       = 112'hC1146E6320696E206E6962682066;
        inPKT[21]       = 112'hC1156163696C6973697320636F6E;
        inPKT[22]       = 112'hC11676616C6C69732E2053656420;
        inPKT[23]       = 112'hC117636F6E6775652068656E6472;
        inPKT[24]       = 112'hC1186572697420696163756C6973;
        inPKT[25]       = 112'hC1192E20566976616D7573207665;
        inPKT[26]       = 112'hC11A686963756C61206C75637475;
        inPKT[27]       = 112'hC11B73206573742C207669746165;
        inPKT[28]       = 112'hC11C207375736369706974206E69;
        inPKT[29]       = 112'hC11D736C20706F72747469746F72;
        inPKT[30]       = 112'hC11E2061632E0D0A0D0A446F6E65;
        inPKT[31]       = 112'hC11F63206D6F6C65737469652073;
        inPKT[32]       = 112'hC120617069656E2069642076756C;
        inPKT[33]       = 112'hC121707574617465207665737469;
        inPKT[34]       = 112'hC12262756C756D2E204E756C6C61;
        inPKT[35]       = 112'hC12320696E206C6967756C612066;
        inPKT[36]       = 112'hC12472696E67696C6C612C20756C;
        inPKT[37]       = 112'hC1256C616D636F72706572207572;
        inPKT[38]       = 112'hC1266E612065742C20706F727474;
        inPKT[39]       = 112'hC12769746F72206C65637475732E;
        inPKT[40]       = 112'hC128205175697371756520626C61;
        inPKT[41]       = 112'hC1296E646974206575206D617572;
        inPKT[42]       = 112'hC12A69732061632068656E647265;
        inPKT[43]       = 112'hC12B7269742E204E756C6C612076;
        inPKT[44]       = 112'hC12C656E656E617469732C206D65;
        inPKT[45]       = 112'hC12D747573206574206C75637475;
        inPKT[46]       = 112'hC12E73206672696E67696C6C612C;
        inPKT[47]       = 112'hC12F206E6962682076656C697420;
        inPKT[48]       = 112'hC130756C6C616D636F7270657220;
        inPKT[49]       = 112'hC1316469616D2C20656765742065;
        inPKT[50]       = 112'hC132666669636974757220697073;
        inPKT[51]       = 112'hC133756D20747572706973206174;
        inPKT[52]       = 112'hC134206E6962682E205574206567;
        inPKT[53]       = 112'hC1356574207072657469756D2065;
        inPKT[54]       = 112'hC136726F732C2065676574206469;
        inPKT[55]       = 112'hC1376374756D206C616375732E20;
        inPKT[56]       = 112'hC1384D616563656E617320757420;
        inPKT[57]       = 112'hC139656E696D2065782E2041656E;
        inPKT[58]       = 112'hC13A65616E207669746165207365;
        inPKT[59]       = 112'hC13B6D7065722066656C69732C20;
        inPKT[60]       = 112'hC13C73656420756C747269636965;
        inPKT[61]       = 112'hC13D732072697375732E20446F6E;
        inPKT[62]       = 112'hC13E656320636F6E736563746574;
        inPKT[63]       = 112'hC13F7572206D69206E69736C2C20;
        inPKT[64]       = 112'hC140617420637572737573206970;
        inPKT[65]       = 112'hC14173756D206772617669646120;
        inPKT[66]       = 112'hC142612E2050686173656C6C7573;
        inPKT[67]       = 112'hC1432073697420616D6574206D61;
        inPKT[68]       = 112'hC144676E612076656C2069707375;
        inPKT[69]       = 112'hC1456D206567657374617320706F;
        inPKT[70]       = 112'hC1467274612E20566976616D7573;
        inPKT[71]       = 112'hC147206C756374757320656E696D;
        inPKT[72]       = 112'hC14820656765742074656D706F72;
        inPKT[73]       = 112'hC1492073616769747469732E2041;
        inPKT[74]       = 112'hC14A6C697175616D20626962656E;
        inPKT[75]       = 112'hC14B64756D2073656D206120636F;
        inPKT[76]       = 112'hC14C6E7365637465747572206566;
        inPKT[77]       = 112'hC14D666963697475722E20446F6E;
        inPKT[78]       = 112'hC14E6563207363656C6572697371;
        inPKT[79]       = 112'hC14F756520616C697175616D2063;
        inPKT[80]       = 112'hC15075727375732E204375726162;
        inPKT[81]       = 112'hC151697475722073697420616D65;
        inPKT[82]       = 112'hC1527420626962656E64756D2065;
        inPKT[83]       = 112'hC1536C69742E2053656420646961;
        inPKT[84]       = 112'hC1546D206A7573746F2C20696163;
        inPKT[85]       = 112'hC155756C69732071756973206E75;
        inPKT[86]       = 112'hC1566C6C612076697461652C2061;
        inPKT[87]       = 112'hC1576C697175616D20657569736D;
        inPKT[88]       = 112'hC1586F642066656C69732E0D0A0D;
        inPKT[89]       = 112'hC1590A50726F696E206461706962;
        inPKT[90]       = 112'hC15A75732C206469616D2076756C;
        inPKT[91]       = 112'hC15B707574617465206672696E67;
        inPKT[92]       = 112'hC15C696C6C61206D616C65737561;
        inPKT[93]       = 112'hC15D64612C206A7573746F207075;
        inPKT[94]       = 112'hC15E72757320636F6D6D6F646F20;
        inPKT[95]       = 112'hC15F646F6C6F722C207574206469;
        inPKT[96]       = 112'hC1606374756D2065726174206E75;
        inPKT[97]       = 112'hC1616E632072757472756D207572;
        inPKT[98]       = 112'hC1626E612E204E756C6C61206772;
        inPKT[99]       = 112'hC16361766964612075726E612076;
        inPKT[100]      = 112'hC1646974616520696D7065726469;
        inPKT[101]      = 112'hC1656574206C616F726565742E20;
        inPKT[102]      = 112'hC16650656C6C656E746573717565;
        inPKT[103]      = 112'hC1672072686F6E63757320626962;
        inPKT[104]      = 112'hC168656E64756D206E6962682C20;
        inPKT[105]      = 112'hC1696964206D6F6C6C6973206469;
        inPKT[106]      = 112'hC16A616D20737573636970697420;
        inPKT[107]      = 112'hC16B61632E2050656C6C656E7465;
        inPKT[108]      = 112'hC16C737175652076656C20696163;
        inPKT[109]      = 112'hC16D756C6973206475692E204D6F;
        inPKT[110]      = 112'hC16E72626920617420616C697175;
        inPKT[111]      = 112'hC16F6574206D617373612E205072;
        inPKT[112]      = 112'hC1706F696E207669746165206F72;
        inPKT[113]      = 112'hC1716E617265206F64696F2C2065;
        inPKT[114]      = 112'hC172752076756C70757461746520;
        inPKT[115]      = 112'hC173697073756D2E2050726F696E;
        inPKT[116]      = 112'hC174206C6F626F727469732C2073;
        inPKT[117]      = 112'hC175656D206E656320657569736D;
        inPKT[118]      = 112'hC1766F642074696E636964756E74;
        inPKT[119]      = 112'hC1772C206175677565206D617572;
        inPKT[120]      = 112'hC1786973207363656C6572697371;
        inPKT[121]      = 112'hC1797565206D61676E612C206574;
        inPKT[122]      = 112'hC17A20706F7375657265206D6920;
        inPKT[123]      = 112'hC17B6E69736C206E6563206E6973;
        inPKT[124]      = 112'hC17C692E20467573636520656C69;
        inPKT[125]      = 112'hC17D74206E657175652C20766172;
        inPKT[126]      = 112'hC17E697573206574206672696E67;
        inPKT[127]      = 112'hC17F696C6C612076697461652C20;
        inPKT[128]      = 112'hC1807661726975732076656C206E;
        inPKT[129]      = 112'hC181657175652E204E756C6C6120;
        inPKT[130]      = 112'hC18265742074656D707573206A75;
        inPKT[131]      = 112'hC18373746F2E204D6F7262692075;
        inPKT[132]      = 112'hC1846C6C616D636F727065722073;
        inPKT[133]      = 112'hC1857573636970697420636F6E67;
        inPKT[134]      = 112'hC18675652E2053656420656C6569;
        inPKT[135]      = 112'hC18766656E64206F64696F206163;
        inPKT[136]      = 112'hC188207375736369706974206469;
        inPKT[137]      = 112'hC189676E697373696D2E20517569;
        inPKT[138]      = 112'hC18A7371756520616E746520656E;
        inPKT[139]      = 112'hC18B696D2C20626C616E64697420;
        inPKT[140]      = 112'hC18C696E20636F6E736571756174;
        inPKT[141]      = 112'hC18D2061632C20696E7465726475;
        inPKT[142]      = 112'hC18E6D2076697461652070757275;
        inPKT[143]      = 112'hC18F732E204D6175726973206575;
        inPKT[144]      = 112'hC19069736D6F6420706F73756572;
        inPKT[145]      = 112'hC19165206C65637475732E205669;
        inPKT[146]      = 112'hC19276616D757320696E74657264;
        inPKT[147]      = 112'hC193756D207175616D2065752073;
        inPKT[148]      = 112'hC194656D70657220666175636962;
        inPKT[149]      = 112'hC19575732E0D0A0D0A496E206D6F;
        inPKT[150]      = 112'hC1966C6573746965206E756C6C61;
        inPKT[151]      = 112'hC19720616E74652C20616320696E;
        inPKT[152]      = 112'hC19874657264756D206D61676E61;
        inPKT[153]      = 112'hC19920636F6E64696D656E74756D;
        inPKT[154]      = 112'hC19A20636F6E64696D656E74756D;
        inPKT[155]      = 112'hC19B2E204475697320756C747269;
        inPKT[156]      = 112'hC19C6369657320736F64616C6573;
        inPKT[157]      = 112'hC19D206E756C6C612C2073697420;
        inPKT[158]      = 112'hC19E616D657420756C6C616D636F;
        inPKT[159]      = 112'hC19F72706572206F64696F207072;
        inPKT[160]      = 112'hC1A0657469756D206E65632E2046;
        inPKT[161]      = 112'hC1A1757363652073656420726973;
        inPKT[162]      = 112'hC1A275732070656C6C656E746573;
        inPKT[163]      = 112'hC1A37175652C20636F6E76616C6C;
        inPKT[164]      = 112'hC1A469732073656D20656765742C;
        inPKT[165]      = 112'hC1A52068656E6472657269742065;
        inPKT[166]      = 112'hC1A67261742E204D6F7262692073;
        inPKT[167]      = 112'hC1A76F64616C6573207665686963;
        inPKT[168]      = 112'hC1A8756C61206C6F626F72746973;
        inPKT[169]      = 112'hC1A92E2041656E65616E20612074;
        inPKT[170]      = 112'hC1AA6F72746F7220637572737573;
        inPKT[171]      = 112'hC1AB2C207363656C657269737175;
        inPKT[172]      = 112'hC1AC65206C6967756C6120706F72;
        inPKT[173]      = 112'hC1AD747469746F722C2065676573;
        inPKT[174]      = 112'hC1AE7461732065726F732E204475;
        inPKT[175]      = 112'hC1AF69732074696E636964756E74;
        inPKT[176]      = 112'hC1B020746F72746F722069642070;
        inPKT[177]      = 112'hC1B16F7375657265206772617669;
        inPKT[178]      = 112'hC1B264612E20496E20636F6E7661;
        inPKT[179]      = 112'hC1B36C6C6973206D692069642069;
        inPKT[180]      = 112'hC1B47073756D206D616C65737561;
        inPKT[181]      = 112'hC1B564612C207574206469637475;
        inPKT[182]      = 112'hC1B66D2065726F7320696D706572;
        inPKT[183]      = 112'hC1B7646965742E2050726F696E20;
        inPKT[184]      = 112'hC1B8756C6C616D636F727065722C;
        inPKT[185]      = 112'hC1B9206D61757269732069642076;
        inPKT[186]      = 112'hC1BA617269757320636F6E677565;
        inPKT[187]      = 112'hC1BB2C2065726F73207361706965;
        inPKT[188]      = 112'hC1BC6E2072686F6E637573206D69;
        inPKT[189]      = 112'hC1BD2C20617420617563746F7220;
        inPKT[190]      = 112'hC1BE6E657175652061726375206C;
        inPKT[191]      = 112'hC1BF616F72656574206469616D2E;
        inPKT[192]      = 112'hC1C00D0A0D0A467573636520706F;
        inPKT[193]      = 112'hC1C172747469746F72206C696265;
        inPKT[194]      = 112'hC1C2726F20617263752C206C6163;
        inPKT[195]      = 112'hC1C3696E69612068656E64726572;
        inPKT[196]      = 112'hC1C46974206469616D20636F6E76;
        inPKT[197]      = 112'hC1C5616C6C6973207365642E2050;
        inPKT[198]      = 112'hC1C6686173656C6C7573206E6F6E;
        inPKT[199]      = 112'hC1C7207475727069732070686172;
        inPKT[200]      = 112'hC1C8657472612C20756C6C616D63;
        inPKT[201]      = 112'hC1C96F72706572206E6571756520;
        inPKT[202]      = 112'hC1CA76656C2C20736F6C6C696369;
        inPKT[203]      = 112'hC1CB747564696E2076656C69742E;
        inPKT[204]      = 112'hC1CC2050656C6C656E7465737175;
        inPKT[205]      = 112'hC1CD65206861626974616E74206D;
        inPKT[206]      = 112'hC1CE6F7262692074726973746971;
        inPKT[207]      = 112'hC1CF75652073656E656374757320;
        inPKT[208]      = 112'hC1D06574206E6574757320657420;
        inPKT[209]      = 112'hC1D16D616C657375616461206661;
        inPKT[210]      = 112'hC1D26D6573206163207475727069;
        inPKT[211]      = 112'hC1D37320656765737461732E204E;
        inPKT[212]      = 112'hC1D4616D206E6563207361706965;
        inPKT[213]      = 112'hC1D56E206D6F6C65737469652C20;
        inPKT[214]      = 112'hC1D664696374756D206D61737361;
        inPKT[215]      = 112'hC1D720656765742C206567657374;
        inPKT[216]      = 112'hC1D86173206F64696F2E20457469;
        inPKT[217]      = 112'hC1D9616D20617263752073617069;
        inPKT[218]      = 112'hC1DA656E2C207072657469756D20;
        inPKT[219]      = 112'hC1DB61206D6F6C6C697320612C20;
        inPKT[220]      = 112'hC1DC76756C707574617465206E6F;
        inPKT[221]      = 112'hC1DD6E20657261742E2055742076;
        inPKT[222]      = 112'hC1DE69746165206E696268206C6F;
        inPKT[223]      = 112'hC1DF626F72746973206C65637475;
        inPKT[224]      = 112'hC1E0732066617563696275732070;
        inPKT[225]      = 112'hC1E16F7274612065752073697420;
        inPKT[226]      = 112'hC1E2616D6574206E69736C2E204D;
        inPKT[227]      = 112'hC1E36F72626920706F7274746974;
        inPKT[228]      = 112'hC1E46F722076656C697420657520;
        inPKT[229]      = 112'hC1E5646F6C6F72206C616F726565;
        inPKT[230]      = 112'hC1E6742C2073697420616D657420;
        inPKT[231]      = 112'hC1E7696D7065726469657420656E;
        inPKT[232]      = 112'hC1E8696D20736F64616C65732E20;
        inPKT[233]      = 112'hC1E94E756C6C616D20756C6C616D;
        inPKT[234]      = 112'hC1EA636F72706572207475727069;
        inPKT[235]      = 112'hC1EB732061742070656C6C656E74;
        inPKT[236]      = 112'hC1EC657371756520766172697573;
        inPKT[237]      = 112'hC1ED2E20566976616D7573206575;
        inPKT[238]      = 112'hC1EE20696D70657264696574206E;
        inPKT[239]      = 112'hC1EF657175652E20536564207175;
        inPKT[240]      = 112'hC1F0697320617563746F7220616E;
        inPKT[241]      = 112'hC1F174652E204D61757269732073;
        inPKT[242]      = 112'hC1F2656D70657220697073756D20;
        inPKT[243]      = 112'hC1F37365642064756920706F7375;
        inPKT[244]      = 112'hC1F46572652C20617420616C6971;
        inPKT[245]      = 112'hC1F575616D206D6574757320656C;
        inPKT[246]      = 112'hC1F6656966656E642E204E756C6C;
        inPKT[247]      = 112'hC1F7616D20747269737469717565;
        inPKT[248]      = 112'hC1F820656C656966656E64206572;
        inPKT[249]      = 112'hC1F96F732C206567657420666572;
        inPKT[250]      = 112'hC1FA6D656E74756D20697073756D;
        inPKT[251]      = 112'hC1FB20656C656D656E74756D206E;
        inPKT[252]      = 112'hC1FC65632E0D0A0D0A50656C6C65;
        inPKT[253]      = 112'hC1FD6E7465737175652068656E64;
        inPKT[254]      = 112'hC1FE726572697420626962656E64;
        inPKT[255]      = 112'hC1FF756D206C6967756C612C2065;
        inPKT[256]      = 112'hC1007420736F64616C6573206D61;
        inPKT[257]      = 112'hC101676E61206461706962757320;
        inPKT[258]      = 112'hC102696E2E20496E20616C697175;
        inPKT[259]      = 112'hC103657420746F72746F72206567;
        inPKT[260]      = 112'hC104657420636F6E736563746574;
        inPKT[261]      = 112'hC105757220636F6E736563746574;
        inPKT[262]      = 112'hC10675722E205175697371756520;
        inPKT[263]      = 112'hC107747269737469717565207269;
        inPKT[264]      = 112'hC10873757320657261742C206574;
        inPKT[265]      = 112'hC10920616C697175657420656C69;
        inPKT[266]      = 112'hC10A7420616C6971756574206575;
        inPKT[267]      = 112'hC10B2E20496E7465676572206E6F;
        inPKT[268]      = 112'hC10C6E206D61676E6120696E2066;
        inPKT[269]      = 112'hC10D656C697320706F7274746974;
        inPKT[270]      = 112'hC10E6F722073616769747469732E;
        inPKT[271]      = 112'hC10F205175697371756520766976;
        inPKT[272]      = 112'hC11065727261206F726369206163;
        inPKT[273]      = 112'hC1112072757472756D206C616F72;
        inPKT[274]      = 112'hC1126565742E2041656E65616E20;
        inPKT[275]      = 112'hC113636F6E76616C6C6973206469;
        inPKT[276]      = 112'hC1146374756D207475727069732C;
        inPKT[277]      = 112'hC1152065742066696E6962757320;
        inPKT[278]      = 112'hC11673617069656E20636F6E6775;
        inPKT[279]      = 112'hC1176520696E2E20536564206120;
        inPKT[280]      = 112'hC11865726174206F726E6172652C;
        inPKT[281]      = 112'hC119206D6F6C6C6973206E69736C;
        inPKT[282]      = 112'hC11A2061632C206469676E697373;
        inPKT[283]      = 112'hC11B696D206E657175652E205175;
        inPKT[284]      = 112'hC11C6973717565206D616C657375;
        inPKT[285]      = 112'hC11D61646120706F737565726520;
        inPKT[286]      = 112'hC11E74757270697320657520756C;
        inPKT[287]      = 112'hC11F6C616D636F727065722E2044;
        inPKT[288]      = 112'hC1206F6E65632076697665727261;
        inPKT[289]      = 112'hC12120626962656E64756D206E75;
        inPKT[290]      = 112'hC1226E632C2064696374756D2069;
        inPKT[291]      = 112'hC1236D70657264696574206E6571;
        inPKT[292]      = 112'hC1247565206D6178696D75732069;
        inPKT[293]      = 112'hC1256E2E20446F6E656320757420;
        inPKT[294]      = 112'hC126756C74726963657320646F6C;
        inPKT[295]      = 112'hC1276F722E20566976616D757320;
        inPKT[296]      = 112'hC128736564206175677565207072;
        inPKT[297]      = 112'hC129657469756D2C20766F6C7574;
        inPKT[298]      = 112'hC12A70617420657261742061632C;
        inPKT[299]      = 112'hC12B20706F727461206469616D2E;
        inPKT[300]      = 112'hC12C204D617572697320696E2070;
        inPKT[301]      = 112'hC12D7572757320756C7472696369;
        inPKT[302]      = 112'hC12E65732C207375736369706974;
        inPKT[303]      = 112'hC12F206469616D207365642C2074;
        inPKT[304]      = 112'hC130696E636964756E7420656E69;
        inPKT[305]      = 112'hC1316D2E20446F6E656320717569;
        inPKT[306]      = 112'hC1327320706F7375657265206E69;
        inPKT[307]      = 112'hC13362682E20496E206861632068;
        inPKT[308]      = 112'hC134616269746173736520706C61;
        inPKT[309]      = 112'hC1357465612064696374756D7374;
        inPKT[310]      = 112'hC1362E0D0A0D0A4D6F726269206F;
        inPKT[311]      = 112'hC137726E617265206A7573746F20;
        inPKT[312]      = 112'hC1386174207175616D2066617563;
        inPKT[313]      = 112'hC139696275732C2073697420616D;
        inPKT[314]      = 112'hC13A6574206D6F6C657374696520;
        inPKT[315]      = 112'hC13B6C656F206375727375732E20;
        inPKT[316]      = 112'hC13C4D6175726973206C616F7265;
        inPKT[317]      = 112'hC13D657420616E74652061206D65;
        inPKT[318]      = 112'hC13E747573206566666963697475;
        inPKT[319]      = 112'hC13F72207661726975732E205365;
        inPKT[320]      = 112'hC140642076656C206F7263692073;
        inPKT[321]      = 112'hC14161676974746973206E756E63;
        inPKT[322]      = 112'hC14220626C616E64697420636F6E;
        inPKT[323]      = 112'hC1437365717561742E2050726165;
        inPKT[324]      = 112'hC14473656E74206D616C65737561;
        inPKT[325]      = 112'hC1456461206E6571756520717569;
        inPKT[326]      = 112'hC146732064696374756D20646967;
        inPKT[327]      = 112'hC1476E697373696D2E20446F6E65;
        inPKT[328]      = 112'hC1486320666163696C6973697320;
        inPKT[329]      = 112'hC14973697420616D65742076656C;
        inPKT[330]      = 112'hC14A6974206575206C6F626F7274;
        inPKT[331]      = 112'hC14B69732E204E756C6C616D2062;
        inPKT[332]      = 112'hC14C6C616E64697420656C656D65;
        inPKT[333]      = 112'hC14D6E74756D206D61757269732C;
        inPKT[334]      = 112'hC14E20766974616520656C656D65;
        inPKT[335]      = 112'hC14F6E74756D20646F6C6F722068;
        inPKT[336]      = 112'hC150656E64726572697420766974;
        inPKT[337]      = 112'hC15161652E204675736365206D6F;
        inPKT[338]      = 112'hC1526C65737469652C20656C6974;
        inPKT[339]      = 112'hC15320757420616C697175657420;
        inPKT[340]      = 112'hC154766F6C75747061742C206E65;
        inPKT[341]      = 112'hC1557175652076656C6974207072;
        inPKT[342]      = 112'hC156657469756D2061756775652C;
        inPKT[343]      = 112'hC157206672696E67696C6C612063;
        inPKT[344]      = 112'hC1586F6E64696D656E74756D206A;
        inPKT[345]      = 112'hC1597573746F2073617069656E20;
        inPKT[346]      = 112'hC15A61206A7573746F2E20506861;
        inPKT[347]      = 112'hC15B73656C6C7573207175697320;
        inPKT[348]      = 112'hC15C617563746F72206C6F72656D;
        inPKT[349]      = 112'hC15D2C20696E20616C697175616D;
        inPKT[350]      = 112'hC15E206E756E632E20557420656C;
        inPKT[351]      = 112'hC15F656966656E6420616E746520;
        inPKT[352]      = 112'hC1606574206E697369206D6F6C65;
        inPKT[353]      = 112'hC1617374696520636F6E76616C6C;
        inPKT[354]      = 112'hC16269732069642065742073656D;
        inPKT[355]      = 112'hC1632E2053656420616320626962;
        inPKT[356]      = 112'hC164656E64756D20617263752E20;
        inPKT[357]      = 112'hC165467573636520766573746962;
        inPKT[358]      = 112'hC166756C756D206E756E63206567;
        inPKT[359]      = 112'hC16765742074656C6C7573206665;
        inPKT[360]      = 112'hC168726D656E74756D2C206E6563;
        inPKT[361]      = 112'hC1692072686F6E637573206D6173;
        inPKT[362]      = 112'hC16A736120636F6D6D6F646F2E20;
        inPKT[363]      = 112'hC16B4D616563656E617320696420;
        inPKT[364]      = 112'hC16C6E756E63206E6F6E20657820;
        inPKT[365]      = 112'hC16D766573746962756C756D206F;
        inPKT[366]      = 112'hC16E726E617265207574206E6563;
        inPKT[367]      = 112'hC16F2065726F732E20416C697175;
        inPKT[368]      = 112'hC170616D20656666696369747572;
        inPKT[369]      = 112'hC17120636F6D6D6F646F20646961;
        inPKT[370]      = 112'hC1726D206964206C6F626F727469;
        inPKT[371]      = 112'hC173732E20536564206163207465;
        inPKT[372]      = 112'hC1746D706F72206C65637475732E;
        inPKT[373]      = 112'hC175204E756E6320656C656D656E;
        inPKT[374]      = 112'hC17674756D207574206C65637475;
        inPKT[375]      = 112'hC177732061632074696E63696475;
        inPKT[376]      = 112'hC1786E742E20557420696163756C;
        inPKT[377]      = 112'hC1796973206E756C6C6120717569;
        inPKT[378]      = 112'hC17A7320657820656C656D656E74;
        inPKT[379]      = 112'hC17B756D2C20616C697175657420;
        inPKT[380]      = 112'hC17C73656D706572206D61676E61;
        inPKT[381]      = 112'hC17D20656C656966656E642E0D0A;
        inPKT[382]      = 112'hC17E0D0A43757261626974757220;
        inPKT[383]      = 112'hC17F746F72746F72206E69736C2C;
        inPKT[384]      = 112'hC18020756C747269636965732069;
        inPKT[385]      = 112'hC1816E206E657175652061632C20;
        inPKT[386]      = 112'hC182616363756D73616E20636F6E;
        inPKT[387]      = 112'hC183736571756174206D65747573;
        inPKT[388]      = 112'hC1842E204D616563656E6173206D;
        inPKT[389]      = 112'hC185617373612073617069656E2C;
        inPKT[390]      = 112'hC186206D617474697320696E2076;
        inPKT[391]      = 112'hC187656E656E6174697320736974;
        inPKT[392]      = 112'hC18820616D65742C20617563746F;
        inPKT[393]      = 112'hC189722073697420616D65742065;
        inPKT[394]      = 112'hC18A6E696D2E204E756E63207669;
        inPKT[395]      = 112'hC18B746165206D6574757320636F;
        inPKT[396]      = 112'hC18C6D6D6F646F2C206D61747469;
        inPKT[397]      = 112'hC18D73206D617373612073697420;
        inPKT[398]      = 112'hC18E616D65742C20766172697573;
        inPKT[399]      = 112'hC18F206C6F72656D2E204E756E63;
        inPKT[400]      = 112'hC19020696E20656C697420656C69;
        inPKT[401]      = 112'hC191742E204E756E63206F726E61;
        inPKT[402]      = 112'hC192726520636F6E736563746574;
        inPKT[403]      = 112'hC1937572206D61676E612C207369;
        inPKT[404]      = 112'hC1947420616D657420706F727474;
        inPKT[405]      = 112'hC19569746F722061726375207268;
        inPKT[406]      = 112'hC1966F6E6375732065752E205375;
        inPKT[407]      = 112'hC1977370656E6469737365207363;
        inPKT[408]      = 112'hC198656C6572697371756520756C;
        inPKT[409]      = 112'hC199747269636965732065782061;
        inPKT[410]      = 112'hC19A20616C697175616D2E205375;
        inPKT[411]      = 112'hC19B7370656E6469737365207275;
        inPKT[412]      = 112'hC19C7472756D20736F6C6C696369;
        inPKT[413]      = 112'hC19D747564696E206E756E632C20;
        inPKT[414]      = 112'hC19E6E6F6E20636F6E76616C6C69;
        inPKT[415]      = 112'hC19F7320747572706973206C616F;
        inPKT[416]      = 112'hC1A0726565742073697420616D65;
        inPKT[417]      = 112'hC1A1742E2041656E65616E206120;
        inPKT[418]      = 112'hC1A266696E69627573206D617572;
        inPKT[419]      = 112'hC1A369732C207175697320637572;
        inPKT[420]      = 112'hC1A4737573206E756E632E20496E;
        inPKT[421]      = 112'hC1A5206665756769617420647569;
        inPKT[422]      = 112'hC1A62076656C2075726E61207365;
        inPKT[423]      = 112'hC1A76D7065722066617563696275;
        inPKT[424]      = 112'hC1A8732E204D617572697320756C;
        inPKT[425]      = 112'hC1A9747269636965732061742074;
        inPKT[426]      = 112'hC1AA757270697320656765742070;
        inPKT[427]      = 112'hC1AB656C6C656E7465737175652E;
        inPKT[428]      = 112'hC1AC205072616573656E74207369;
        inPKT[429]      = 112'hC1AD7420616D6574206C6967756C;
        inPKT[430]      = 112'hC1AE6120636F6E76616C6C69732C;
        inPKT[431]      = 112'hC1AF20656C656D656E74756D206E;
        inPKT[432]      = 112'hC1B0756C6C6120756C6C616D636F;
        inPKT[433]      = 112'hC1B1727065722C20616C69717561;
        inPKT[434]      = 112'hC1B26D2075726E612E2045746961;
        inPKT[435]      = 112'hC1B36D207175616D20656C69742C;
        inPKT[436]      = 112'hC1B420706F737565726520757420;
        inPKT[437]      = 112'hC1B57175616D20656765742C2066;
        inPKT[438]      = 112'hC1B6696E6962757320736F6C6C69;
        inPKT[439]      = 112'hC1B76369747564696E206E756C6C;
        inPKT[440]      = 112'hC1B8612E20496E20737573636970;
        inPKT[441]      = 112'hC1B9697420656E696D2065742065;
        inPKT[442]      = 112'hC1BA726F732066696E696275732C;
        inPKT[443]      = 112'hC1BB207574207363656C65726973;
        inPKT[444]      = 112'hC1BC7175652074656C6C75732066;
        inPKT[445]      = 112'hC1BD6575676961742E2043757261;
        inPKT[446]      = 112'hC1BE6269747572206E6F6E206D61;
        inPKT[447]      = 112'hC1BF737361207661726975732064;
        inPKT[448]      = 112'hC1C06F6C6F722067726176696461;
        inPKT[449]      = 112'hC1C120656C656D656E74756D2071;
        inPKT[450]      = 112'hC1C27569732075742066656C6973;
        inPKT[451]      = 112'hC1C32E2050686173656C6C757320;
        inPKT[452]      = 112'hC1C4657569736D6F642069707375;
        inPKT[453]      = 112'hC1C56D20656765742076656C6974;
        inPKT[454]      = 112'hC1C6206C6F626F727469732C2065;
        inPKT[455]      = 112'hC1C767657420706F727461206D61;
        inPKT[456]      = 112'hC1C8757269732074656D7075732E;
        inPKT[457]      = 112'hC1C92053656420696D7065726469;
        inPKT[458]      = 112'hC1CA657420766F6C757470617420;
        inPKT[459]      = 112'hC1CB74656C6C7573206575207469;
        inPKT[460]      = 112'hC1CC6E636964756E742E0D0A0D0A;
        inPKT[461]      = 112'hC1CD55742076656C206D69206174;
        inPKT[462]      = 112'hC1CE206D65747573206672696E67;
        inPKT[463]      = 112'hC1CF696C6C612067726176696461;
        inPKT[464]      = 112'hC1D02E205072616573656E742065;
        inPKT[465]      = 112'hC1D1726F73206E6962682C206375;
        inPKT[466]      = 112'hC1D2727375732065676573746173;
        inPKT[467]      = 112'hC1D32074696E636964756E742073;
        inPKT[468]      = 112'hC1D46F64616C65732C207363656C;
        inPKT[469]      = 112'hC1D565726973717565206E656320;
        inPKT[470]      = 112'hC1D666656C69732E20496E746567;
        inPKT[471]      = 112'hC1D7657220696D70657264696574;
        inPKT[472]      = 112'hC1D8206D616C657375616461206E;
        inPKT[473]      = 112'hC1D969736C20616C697175657420;
        inPKT[474]      = 112'hC1DA76656E656E617469732E2049;
        inPKT[475]      = 112'hC1DB6E7465676572207365642070;
        inPKT[476]      = 112'hC1DC6F72747469746F7220697073;
        inPKT[477]      = 112'hC1DD756D2E20496E746567657220;
        inPKT[478]      = 112'hC1DE636F6D6D6F646F2066657567;
        inPKT[479]      = 112'hC1DF69617420746F72746F722C20;
        inPKT[480]      = 112'hC1E06575206C6F626F7274697320;
        inPKT[481]      = 112'hC1E1617567756520656C656D656E;
        inPKT[482]      = 112'hC1E274756D2073697420616D6574;
        inPKT[483]      = 112'hC1E32E20446F6E65632076657374;
        inPKT[484]      = 112'hC1E46962756C756D206C6967756C;
        inPKT[485]      = 112'hC1E5612061756775652C20657420;
        inPKT[486]      = 112'hC1E666696E696275732061726375;
        inPKT[487]      = 112'hC1E720706F72746120696E2E204E;
        inPKT[488]      = 112'hC1E8756C6C612073656D2074656C;
        inPKT[489]      = 112'hC1E96C75732C20756C6C616D636F;
        inPKT[490]      = 112'hC1EA727065722061742063757273;
        inPKT[491]      = 112'hC1EB757320612C20706F72746120;
        inPKT[492]      = 112'hC1EC73697420616D6574206D6167;
        inPKT[493]      = 112'hC1ED6E612E204E756E6320766974;
        inPKT[494]      = 112'hC1EE616520696D70657264696574;
        inPKT[495]      = 112'hC1EF2070757275732C206E656320;
        inPKT[496]      = 112'hC1F0736F6C6C696369747564696E;
        inPKT[497]      = 112'hC1F12074656C6C75732E20416C69;
        inPKT[498]      = 112'hC1F27175616D206572617420766F;
        inPKT[499]      = 112'hC1F36C75747061742E2053656420;
        inPKT[500]      = 112'hC1F46964206D61676E6120636F6D;
        inPKT[501]      = 112'hC1F56D6F646F2C206C7563747573;
        inPKT[502]      = 112'hC1F62076656C697420717569732C;
        inPKT[503]      = 112'hC1F720657569736D6F6420656E69;
        inPKT[504]      = 112'hC1F86D2E20496E7465676572206D;
        inPKT[505]      = 112'hC1F9617474697320736F64616C65;
        inPKT[506]      = 112'hC1FA73206665726D656E74756D2E;
        inPKT[507]      = 112'hC1FB205175697371756520736564;
        inPKT[508]      = 112'hC1FC206672696E67696C6C61206C;
        inPKT[509]      = 112'hC1FD6F72656D2E20437261732076;
        inPKT[510]      = 112'hC1FE65686963756C612074656D70;
        inPKT[511]      = 112'hC1FF75732073617069656E207574;
        inPKT[512]      = 112'hC10020636F6E6775652E20447569;
        inPKT[513]      = 112'hC101732073617069656E20656E69;
        inPKT[514]      = 112'hC1026D2C20706F727461206E6563;
        inPKT[515]      = 112'hC103206C656F2069642C20656666;
        inPKT[516]      = 112'hC10469636974757220706F737565;
        inPKT[517]      = 112'hC1057265206C696265726F2E204E;
        inPKT[518]      = 112'hC106756C6C616D2061632074656D;
        inPKT[519]      = 112'hC107706F72206D657475732E2053;
        inPKT[520]      = 112'hC10865642076656C207475727069;
        inPKT[521]      = 112'hC1097320666575676961742C2069;
        inPKT[522]      = 112'hC10A6163756C6973206175677565;
        inPKT[523]      = 112'hC10B20717569732C2074696E6369;
        inPKT[524]      = 112'hC10C64756E74207475727069732E;
        inPKT[525]      = 112'hC10D0D0A0D0A566976616D757320;
        inPKT[526]      = 112'hC10E706F737565726520706F7274;
        inPKT[527]      = 112'hC10F7469746F722061756775652C;
        inPKT[528]      = 112'hC110207661726975732061636375;
        inPKT[529]      = 112'hC1116D73616E20656C6974207675;
        inPKT[530]      = 112'hC1126C7075746174652065676574;
        inPKT[531]      = 112'hC1132E2051756973717565207365;
        inPKT[532]      = 112'hC11464206D616C65737561646120;
        inPKT[533]      = 112'hC1156E69736C2E20496E74657264;
        inPKT[534]      = 112'hC116756D206574206D616C657375;
        inPKT[535]      = 112'hC1176164612066616D6573206163;
        inPKT[536]      = 112'hC11820616E746520697073756D20;
        inPKT[537]      = 112'hC1197072696D697320696E206661;
        inPKT[538]      = 112'hC11A7563696275732E204E756E63;
        inPKT[539]      = 112'hC11B20747572706973206469616D;
        inPKT[540]      = 112'hC11C2C2073757363697069742061;
        inPKT[541]      = 112'hC11D632065726F732076656C2C20;
        inPKT[542]      = 112'hC11E74656D7075732076656E656E;
        inPKT[543]      = 112'hC11F6174697320697073756D2E20;
        inPKT[544]      = 112'hC12044756973206C756374757320;
        inPKT[545]      = 112'hC12172686F6E637573206D617373;
        inPKT[546]      = 112'hC122612E20467573636520757420;
        inPKT[547]      = 112'hC1236C6163696E69612074757270;
        inPKT[548]      = 112'hC12469732E20566976616D757320;
        inPKT[549]      = 112'hC12572757472756D2074656C6C75;
        inPKT[550]      = 112'hC126732061756775652C20617420;
        inPKT[551]      = 112'hC1276F726E617265206E69736C20;
        inPKT[552]      = 112'hC128666163696C69736973206574;
        inPKT[553]      = 112'hC1292E204E756E6320736564206E;
        inPKT[554]      = 112'hC12A6973692072697375732E2049;
        inPKT[555]      = 112'hC12B6E746567657220656C656D65;
        inPKT[556]      = 112'hC12C6E74756D206D617572697320;
        inPKT[557]      = 112'hC12D7175616D2C20757420766568;
        inPKT[558]      = 112'hC12E6963756C61206D6175726973;
        inPKT[559]      = 112'hC12F20636F6E6775652065752E0D;
        inPKT[560]      = 112'hC1300A0D0A467573636520612074;
        inPKT[561]      = 112'hC131656C6C75732073697420616D;
        inPKT[562]      = 112'hC13265742065726174206665726D;
        inPKT[563]      = 112'hC133656E74756D207363656C6572;
        inPKT[564]      = 112'hC13469737175652E204375726162;
        inPKT[565]      = 112'hC1356974757220696E2076656C69;
        inPKT[566]      = 112'hC1367420617420656E696D206C61;
        inPKT[567]      = 112'hC13763696E696120766568696375;
        inPKT[568]      = 112'hC1386C61206163206964206A7573;
        inPKT[569]      = 112'hC139746F2E2050726F696E206E6F;
        inPKT[570]      = 112'hC13A6E20646F6C6F722065666669;
        inPKT[571]      = 112'hC13B63697475722C2074696E6369;
        inPKT[572]      = 112'hC13C64756E74206F64696F206575;
        inPKT[573]      = 112'hC13D2C2066617563696275732065;
        inPKT[574]      = 112'hC13E6E696D2E2050656C6C656E74;
        inPKT[575]      = 112'hC13F657371756520646170696275;
        inPKT[576]      = 112'hC14073206F726369206163206C6F;
        inPKT[577]      = 112'hC14172656D20696163756C69732C;
        inPKT[578]      = 112'hC1422073697420616D657420626C;
        inPKT[579]      = 112'hC143616E64697420617263752074;
        inPKT[580]      = 112'hC14472697374697175652E204165;
        inPKT[581]      = 112'hC1456E65616E2074726973746971;
        inPKT[582]      = 112'hC146756520746F72746F72206E65;
        inPKT[583]      = 112'hC14763206A7573746F20616C6971;
        inPKT[584]      = 112'hC14875616D2C20696E2070726574;
        inPKT[585]      = 112'hC14969756D2066656C6973206D6F;
        inPKT[586]      = 112'hC14A6C65737469652E2053656420;
        inPKT[587]      = 112'hC14B65742074656D707573206175;
        inPKT[588]      = 112'hC14C6775652E204E756C6C612066;
        inPKT[589]      = 112'hC14D72696E67696C6C6120656C65;
        inPKT[590]      = 112'hC14E6966656E6420697073756D20;
        inPKT[591]      = 112'hC14F766976657272612063757273;
        inPKT[592]      = 112'hC15075732E20416C697175616D20;
        inPKT[593]      = 112'hC1516D6178696D7573206665726D;
        inPKT[594]      = 112'hC152656E74756D206E6962682061;
        inPKT[595]      = 112'hC1536320616363756D73616E2E20;
        inPKT[596]      = 112'hC1544E756C6C6120666163696C69;
        inPKT[597]      = 112'hC15573692E20566573746962756C;
        inPKT[598]      = 112'hC156756D20666163696C69736973;
        inPKT[599]      = 112'hC157206C656F2065676573746173;
        inPKT[600]      = 112'hC1582073656D206D617474697320;
        inPKT[601]      = 112'hC159636F6E6775652E204D617572;
        inPKT[602]      = 112'hC15A697320766974616520657820;
        inPKT[603]      = 112'hC15B617420726973757320646170;
        inPKT[604]      = 112'hC15C6962757320656C656966656E;
        inPKT[605]      = 112'hC15D642E20496E74656765722075;
        inPKT[606]      = 112'hC15E742065726F7320636F6E6775;
        inPKT[607]      = 112'hC15F652C20706F72747469746F72;
        inPKT[608]      = 112'hC16020616E7465206E6F6E2C2069;
        inPKT[609]      = 112'hC1616E74657264756D20646F6C6F;
        inPKT[610]      = 112'hC162722E0D0A0D0A566573746962;
        inPKT[611]      = 112'hC163756C756D20656C656966656E;
        inPKT[612]      = 112'hC16464206D617572697320657520;
        inPKT[613]      = 112'hC1656E6973692064696374756D20;
        inPKT[614]      = 112'hC166677261766964612E20447569;
        inPKT[615]      = 112'hC16773206D6F6C6C697320646961;
        inPKT[616]      = 112'hC1686D2076656C20656E696D2074;
        inPKT[617]      = 112'hC169656D7075732C207669746165;
        inPKT[618]      = 112'hC16A2064617069627573206D6173;
        inPKT[619]      = 112'hC16B73612073616769747469732E;
        inPKT[620]      = 112'hC16C204E756C6C61207574206175;
        inPKT[621]      = 112'hC16D63746F7220746F72746F722E;
        inPKT[622]      = 112'hC16E204D6F72626920736564206C;
        inPKT[623]      = 112'hC16F6F72656D2075726E612E2046;
        inPKT[624]      = 112'hC17075736365206D61747469732C;
        inPKT[625]      = 112'hC171206D61676E6120616320636F;
        inPKT[626]      = 112'hC1726E64696D656E74756D206665;
        inPKT[627]      = 112'hC17375676961742C206D61737361;
        inPKT[628]      = 112'hC17420647569206D6178696D7573;
        inPKT[629]      = 112'hC175206E756C6C612C2065752061;
        inPKT[630]      = 112'hC1766C6971756574206E65717565;
        inPKT[631]      = 112'hC177206D61757269732061206572;
        inPKT[632]      = 112'hC17861742E205175697371756520;
        inPKT[633]      = 112'hC179617563746F72206573742075;
        inPKT[634]      = 112'hC17A7420696E74657264756D2063;
        inPKT[635]      = 112'hC17B6F6E73656374657475722E20;
        inPKT[636]      = 112'hC17C446F6E656320656765742064;
        inPKT[637]      = 112'hC17D69676E697373696D20746F72;
        inPKT[638]      = 112'hC17E746F722C2068656E64726572;
        inPKT[639]      = 112'hC17F6974206D6174746973206572;
        inPKT[640]      = 112'hC18061742E2050656C6C656E7465;
        inPKT[641]      = 112'hC18173717565206861626974616E;
        inPKT[642]      = 112'hC18274206D6F7262692074726973;
        inPKT[643]      = 112'hC18374697175652073656E656374;
        inPKT[644]      = 112'hC1847573206574206E6574757320;
        inPKT[645]      = 112'hC1856574206D616C657375616461;
        inPKT[646]      = 112'hC1862066616D6573206163207475;
        inPKT[647]      = 112'hC187727069732065676573746173;
        inPKT[648]      = 112'hC1882E2051756973717565206F72;
        inPKT[649]      = 112'hC1896E6172652076617269757320;
        inPKT[650]      = 112'hC18A74656D7075732E0D0A0D0A4D;
        inPKT[651]      = 112'hC18B6F7262692072757472756D20;
        inPKT[652]      = 112'hC18C616E7465206E6962682C2061;
        inPKT[653]      = 112'hC18D2076697665727261206E756C;
        inPKT[654]      = 112'hC18E6C612068656E647265726974;
        inPKT[655]      = 112'hC18F20696E2E2050726F696E2073;
        inPKT[656]      = 112'hC190757363697069742065676573;
        inPKT[657]      = 112'hC19174617320657261742C207574;
        inPKT[658]      = 112'hC19220617563746F72206F726369;
        inPKT[659]      = 112'hC193206D617474697320612E2050;
        inPKT[660]      = 112'hC194656C6C656E74657371756520;
        inPKT[661]      = 112'hC1956C7563747573206672696E67;
        inPKT[662]      = 112'hC196696C6C6120656C6974207574;
        inPKT[663]      = 112'hC197206C6163696E69612E205574;
        inPKT[664]      = 112'hC198206574206D61737361206E75;
        inPKT[665]      = 112'hC1996C6C612E2053656420617420;
        inPKT[666]      = 112'hC19A6672696E67696C6C61206C6F;
        inPKT[667]      = 112'hC19B72656D2E2050726F696E2067;
        inPKT[668]      = 112'hC19C72617669646120616363756D;
        inPKT[669]      = 112'hC19D73616E207269737573207365;
        inPKT[670]      = 112'hC19E6420626962656E64756D2E20;
        inPKT[671]      = 112'hC19F4D616563656E6173206D616C;
        inPKT[672]      = 112'hC1A0657375616461206F64696F20;
        inPKT[673]      = 112'hC1A175742076656C697420657569;
        inPKT[674]      = 112'hC1A2736D6F642064617069627573;
        inPKT[675]      = 112'hC1A32E0D0A0D0A457469616D2063;
        inPKT[676]      = 112'hC1A46F6E677565206D6174746973;
        inPKT[677]      = 112'hC1A520696163756C69732E204D61;
        inPKT[678]      = 112'hC1A6757269732076697461652065;
        inPKT[679]      = 112'hC1A766666963697475722073656D;
        inPKT[680]      = 112'hC1A82E205365642070756C76696E;
        inPKT[681]      = 112'hC1A9617220646F6C6F7220757420;
        inPKT[682]      = 112'hC1AA6D6920657569736D6F642068;
        inPKT[683]      = 112'hC1AB656E6472657269742E204E75;
        inPKT[684]      = 112'hC1AC6C6C616D2061742067726176;
        inPKT[685]      = 112'hC1AD69646120646F6C6F722E204D;
        inPKT[686]      = 112'hC1AE6F726269206C656F20747572;
        inPKT[687]      = 112'hC1AF7069732C20636F6E67756520;
        inPKT[688]      = 112'hC1B06E656320616C697175616D20;
        inPKT[689]      = 112'hC1B175742C20636F6D6D6F646F20;
        inPKT[690]      = 112'hC1B2696E206E756E632E204E756C;
        inPKT[691]      = 112'hC1B36C6120617420666175636962;
        inPKT[692]      = 112'hC1B47573206C656F2C2065752066;
        inPKT[693]      = 112'hC1B5657567696174206C61637573;
        inPKT[694]      = 112'hC1B62E204675736365206E6F6E20;
        inPKT[695]      = 112'hC1B7656765737461732074757270;
        inPKT[696]      = 112'hC1B869732E205175697371756520;
        inPKT[697]      = 112'hC1B9766974616520697073756D20;
        inPKT[698]      = 112'hC1BA6D692E204E756E63206E6F6E;
        inPKT[699]      = 112'hC1BB206F7263692073697420616D;
        inPKT[700]      = 112'hC1BC6574206E6973692076617269;
        inPKT[701]      = 112'hC1BD757320706F72747469746F72;
        inPKT[702]      = 112'hC1BE20696E2076756C7075746174;
        inPKT[703]      = 112'hC1BF6520746F72746F722E204E75;
        inPKT[704]      = 112'hC1C06E6320636F6E76616C6C6973;
        inPKT[705]      = 112'hC1C1206772617669646120646961;
        inPKT[706]      = 112'hC1C26D206120756C747269636965;
        inPKT[707]      = 112'hC1C3732E20517569737175652065;
        inPKT[708]      = 112'hC1C475206A7573746F20636F6E64;
        inPKT[709]      = 112'hC1C5696D656E74756D2C20766172;
        inPKT[710]      = 112'hC1C6697573206469616D2076656C;
        inPKT[711]      = 112'hC1C72C20766573746962756C756D;
        inPKT[712]      = 112'hC1C8206D617373612E0D0A0D0A50;
        inPKT[713]      = 112'hC1C9656C6C656E74657371756520;
        inPKT[714]      = 112'hC1CA70656C6C656E746573717565;
        inPKT[715]      = 112'hC1CB2073617069656E206E657175;
        inPKT[716]      = 112'hC1CC652C20617563746F72206D61;
        inPKT[717]      = 112'hC1CD6C6573756164612065726174;
        inPKT[718]      = 112'hC1CE2068656E647265726974206E;
        inPKT[719]      = 112'hC1CF65632E204E756C6C6120706C;
        inPKT[720]      = 112'hC1D0616365726174206469616D20;
        inPKT[721]      = 112'hC1D168656E647265726974206D61;
        inPKT[722]      = 112'hC1D273736120626962656E64756D;
        inPKT[723]      = 112'hC1D32C2061206D6F6C6573746965;
        inPKT[724]      = 112'hC1D42066656C69732068656E6472;
        inPKT[725]      = 112'hC1D5657269742E204D6175726973;
        inPKT[726]      = 112'hC1D620657569736D6F642076656E;
        inPKT[727]      = 112'hC1D7656E61746973206A7573746F;
        inPKT[728]      = 112'hC1D82C20757420617563746F7220;
        inPKT[729]      = 112'hC1D9656C697420616C6971756574;
        inPKT[730]      = 112'hC1DA2075742E2046757363652061;
        inPKT[731]      = 112'hC1DB6C69717565742C207175616D;
        inPKT[732]      = 112'hC1DC207574206469676E69737369;
        inPKT[733]      = 112'hC1DD6D2068656E6472657269742C;
        inPKT[734]      = 112'hC1DE206D61757269732074757270;
        inPKT[735]      = 112'hC1DF6973206469676E697373696D;
        inPKT[736]      = 112'hC1E020746F72746F722C20656765;
        inPKT[737]      = 112'hC1E1742070656C6C656E74657371;
        inPKT[738]      = 112'hC1E275652076656C6974206F7263;
        inPKT[739]      = 112'hC1E369206E6563207175616D2E20;
        inPKT[740]      = 112'hC1E44E756E632065676573746173;
        inPKT[741]      = 112'hC1E52070656C6C656E7465737175;
        inPKT[742]      = 112'hC1E6652072697375732E20437572;
        inPKT[743]      = 112'hC1E7616269747572207375736369;
        inPKT[744]      = 112'hC1E87069742074656D707573206C;
        inPKT[745]      = 112'hC1E9616375732C20656765742070;
        inPKT[746]      = 112'hC1EA72657469756D20656C697420;
        inPKT[747]      = 112'hC1EB74696E636964756E74206E6F;
        inPKT[748]      = 112'hC1EC6E2E20437261732075726E61;
        inPKT[749]      = 112'hC1ED206C6F72656D2C20706C6163;
        inPKT[750]      = 112'hC1EE6572617420766F6C75747061;
        inPKT[751]      = 112'hC1EF7420696D7065726469657420;
        inPKT[752]      = 112'hC1F073697420616D65742C206567;
        inPKT[753]      = 112'hC1F165737461732076656C206F72;
        inPKT[754]      = 112'hC1F263692E0D0A0D0A50656C6C65;
        inPKT[755]      = 112'hC1F36E74657371756520736F6461;
        inPKT[756]      = 112'hC1F46C6573206665726D656E7475;
        inPKT[757]      = 112'hC1F56D206E69736C2C2061742066;
        inPKT[758]      = 112'hC1F672696E67696C6C6120647569;
        inPKT[759]      = 112'hC1F72073656D706572206665726D;
        inPKT[760]      = 112'hC1F8656E74756D2E204E756C6C61;
        inPKT[761]      = 112'hC1F96D20706C6163657261742076;
        inPKT[762]      = 112'hC1FA656C206D692068656E647265;
        inPKT[763]      = 112'hC1FB72697420656C656D656E7475;
        inPKT[764]      = 112'hC1FC6D2E20457469616D206E6F6E;
        inPKT[765]      = 112'hC1FD20697073756D2065782E204E;
        inPKT[766]      = 112'hC1FE616D206163207363656C6572;
        inPKT[767]      = 112'hC1FF6973717565206E6962682C20;
        inPKT[768]      = 112'hC10076656C20666163696C697369;
        inPKT[769]      = 112'hC10173206D692E20446F6E656320;
        inPKT[770]      = 112'hC10265676573746173206C616F72;
        inPKT[771]      = 112'hC1036565742065726F732C206567;
        inPKT[772]      = 112'hC104657420766F6C757470617420;
        inPKT[773]      = 112'hC1056D657475732E205072616573;
        inPKT[774]      = 112'hC106656E7420616363756D73616E;
        inPKT[775]      = 112'hC10720626962656E64756D206E69;
        inPKT[776]      = 112'hC108736C206E65632076656E656E;
        inPKT[777]      = 112'hC109617469732E20536564207275;
        inPKT[778]      = 112'hC10A7472756D206D692061207375;
        inPKT[779]      = 112'hC10B736369706974207068617265;
        inPKT[780]      = 112'hC10C7472612E2053656420736974;
        inPKT[781]      = 112'hC10D20616D657420696E74657264;
        inPKT[782]      = 112'hC10E756D207475727069732E2041;
        inPKT[783]      = 112'hC10F6C697175616D206575206E69;
        inPKT[784]      = 112'hC110626820746F72746F722E2044;
        inPKT[785]      = 112'hC1116F6E65632066617563696275;
        inPKT[786]      = 112'hC112732064617069627573206E69;
        inPKT[787]      = 112'hC11373692C20736564206C616F72;
        inPKT[788]      = 112'hC114656574206F72636920736365;
        inPKT[789]      = 112'hC1156C6572697371756520696E2E;
        inPKT[790]      = 112'hC1160D0A0D0A4D61757269732069;
        inPKT[791]      = 112'hC1176E2066656C6973206665726D;
        inPKT[792]      = 112'hC118656E74756D2C20636F6E7661;
        inPKT[793]      = 112'hC1196C6C69732061756775652076;
        inPKT[794]      = 112'hC11A656C2C20706F737565726520;
        inPKT[795]      = 112'hC11B6D692E2050656C6C656E7465;
        inPKT[796]      = 112'hC11C73717565207363656C657269;
        inPKT[797]      = 112'hC11D737175652072686F6E637573;
        inPKT[798]      = 112'hC11E206A7573746F2C2065752070;
        inPKT[799]      = 112'hC11F756C76696E617220656E696D;
        inPKT[800]      = 112'hC1202070756C76696E6172207665;
        inPKT[801]      = 112'hC1216C2E204D616563656E617320;
        inPKT[802]      = 112'hC1227068617265747261206C6962;
        inPKT[803]      = 112'hC12365726F206D61676E612C2061;
        inPKT[804]      = 112'hC1246320736F6C6C696369747564;
        inPKT[805]      = 112'hC125696E206C656F206D6F6C6C69;
        inPKT[806]      = 112'hC12673206E6F6E2E204E756C6C61;
        inPKT[807]      = 112'hC12720656C656D656E74756D206F;
        inPKT[808]      = 112'hC128726E61726520656765737461;
        inPKT[809]      = 112'hC129732E20436C61737320617074;
        inPKT[810]      = 112'hC12A656E74207461636974692073;
        inPKT[811]      = 112'hC12B6F63696F737175206164206C;
        inPKT[812]      = 112'hC12C69746F726120746F72717565;
        inPKT[813]      = 112'hC12D6E742070657220636F6E7562;
        inPKT[814]      = 112'hC12E6961206E6F737472612C2070;
        inPKT[815]      = 112'hC12F657220696E636570746F7320;
        inPKT[816]      = 112'hC13068696D656E61656F732E2050;
        inPKT[817]      = 112'hC13172616573656E742061756775;
        inPKT[818]      = 112'hC13265206D61757269732C207268;
        inPKT[819]      = 112'hC1336F6E63757320717569732065;
        inPKT[820]      = 112'hC1347374206E6F6E2C206D6F6C6C;
        inPKT[821]      = 112'hC135697320636F6E76616C6C6973;
        inPKT[822]      = 112'hC1362066656C69732E2053757370;
        inPKT[823]      = 112'hC137656E64697373652066616369;
        inPKT[824]      = 112'hC1386C697369732C206F72636920;
        inPKT[825]      = 112'hC1397669746165206C6163696E69;
        inPKT[826]      = 112'hC13A612074656D706F722C206C65;
        inPKT[827]      = 112'hC13B637475732073617069656E20;
        inPKT[828]      = 112'hC13C6D6174746973207269737573;
        inPKT[829]      = 112'hC13D2C206E6F6E20736167697474;
        inPKT[830]      = 112'hC13E697320656C6974206E657175;
        inPKT[831]      = 112'hC13F652071756973206A7573746F;
        inPKT[832]      = 112'hC1402E20446F6E6563206D616C65;
        inPKT[833]      = 112'hC1417375616461206C6163696E69;
        inPKT[834]      = 112'hC14261206475692E205068617365;
        inPKT[835]      = 112'hC1436C6C75732068656E64726572;
        inPKT[836]      = 112'hC1446974206D6175726973206D61;
        inPKT[837]      = 112'hC145757269732C20736564206672;
        inPKT[838]      = 112'hC146696E67696C6C61206C696265;
        inPKT[839]      = 112'hC147726F206672696E67696C6C61;
        inPKT[840]      = 112'hC14820696E2E2053656420617420;
        inPKT[841]      = 112'hC1496C6967756C6120696E206A75;
        inPKT[842]      = 112'hC14A73746F2066696E6962757320;
        inPKT[843]      = 112'hC14B76756C7075746174652E204E;
        inPKT[844]      = 112'hC14C756E6320637572737573206E;
        inPKT[845]      = 112'hC14D657175652073697420616D65;
        inPKT[846]      = 112'hC14E7420617263752074696E6369;
        inPKT[847]      = 112'hC14F64756E742C20766974616520;
        inPKT[848]      = 112'hC15070686172657472612073656D;
        inPKT[849]      = 112'hC15120706F72747469746F722E20;
        inPKT[850]      = 112'hC152416C697175616D206D617474;
        inPKT[851]      = 112'hC15369732C206A7573746F206E6F;
        inPKT[852]      = 112'hC1546E20657569736D6F6420636F;
        inPKT[853]      = 112'hC1556E76616C6C69732C206E756E;
        inPKT[854]      = 112'hC15663206D6920636F6E73657175;
        inPKT[855]      = 112'hC1576174206573742C206E656320;
        inPKT[856]      = 112'hC158736F6C6C696369747564696E;
        inPKT[857]      = 112'hC159206C65637475732073617069;
        inPKT[858]      = 112'hC15A656E2076656C206F64696F2E;
        inPKT[859]      = 112'hC15B20496E2074656D706F722065;
        inPKT[860]      = 112'hC15C72617420646F6C6F722C2073;
        inPKT[861]      = 112'hC15D6564207665686963756C6120;
        inPKT[862]      = 112'hC15E75726E6120636F6E73657175;
        inPKT[863]      = 112'hC15F6174207365642E0D0A0D0A4E;
        inPKT[864]      = 112'hC160616D2072686F6E6375732069;
        inPKT[865]      = 112'hC16164206D6175726973206E6563;
        inPKT[866]      = 112'hC162206469676E697373696D2E20;
        inPKT[867]      = 112'hC163496E20696D70657264696574;
        inPKT[868]      = 112'hC16420756C747269636573206572;
        inPKT[869]      = 112'hC1656174206E656320736F6C6C69;
        inPKT[870]      = 112'hC1666369747564696E2E20496E74;
        inPKT[871]      = 112'hC167656765722073656420636F6E;
        inPKT[872]      = 112'hC16864696D656E74756D2065726F;
        inPKT[873]      = 112'hC169732E20446F6E656320656765;
        inPKT[874]      = 112'hC16A74206E756E63206964206D61;
        inPKT[875]      = 112'hC16B757269732074726973746971;
        inPKT[876]      = 112'hC16C756520706F72747469746F72;
        inPKT[877]      = 112'hC16D206C616F7265657420766974;
        inPKT[878]      = 112'hC16E6165206D657475732E204E75;
        inPKT[879]      = 112'hC16F6C6C6120666163696C697369;
        inPKT[880]      = 112'hC1702E204E756C6C616D20657520;
        inPKT[881]      = 112'hC1716C616375732061206469616D;
        inPKT[882]      = 112'hC172207472697374697175652065;
        inPKT[883]      = 112'hC173676573746173206E6F6E2069;
        inPKT[884]      = 112'hC1746163756C6973206D65747573;
        inPKT[885]      = 112'hC1752E20416C697175616D20696E;
        inPKT[886]      = 112'hC1762074656D706F722065726174;
        inPKT[887]      = 112'hC1772C20696420636F6E67756520;
        inPKT[888]      = 112'hC1786D617373612E20566976616D;
        inPKT[889]      = 112'hC17975732076656C20746F72746F;
        inPKT[890]      = 112'hC17A72207669746165206E696268;
        inPKT[891]      = 112'hC17B20636F6D6D6F646F206C6F62;
        inPKT[892]      = 112'hC17C6F7274697320717569732061;
        inPKT[893]      = 112'hC17D20697073756D2E2050726F69;
        inPKT[894]      = 112'hC17E6E20766F6C75747061742071;
        inPKT[895]      = 112'hC17F75616D206E6F6E2066656C69;
        inPKT[896]      = 112'hC180732074656D7075732C206964;
        inPKT[897]      = 112'hC18120706F737565726520646F6C;
        inPKT[898]      = 112'hC1826F722074656D706F722E2050;
        inPKT[899]      = 112'hC18372616573656E742076697461;
        inPKT[900]      = 112'hC184652074696E636964756E7420;
        inPKT[901]      = 112'hC18573617069656E2E204D616563;
        inPKT[902]      = 112'hC186656E617320666163696C6973;
        inPKT[903]      = 112'hC1876973206D617474697320616E;
        inPKT[904]      = 112'hC188746520717569732076617269;
        inPKT[905]      = 112'hC18975732E20446F6E6563207065;
        inPKT[906]      = 112'hC18A6C6C656E7465737175652065;
        inPKT[907]      = 112'hC18B726F73206665756769617420;
        inPKT[908]      = 112'hC18C74696E636964756E7420636F;
        inPKT[909]      = 112'hC18D6E64696D656E74756D2E2050;
        inPKT[910]      = 112'hC18E726F696E2066617563696275;
        inPKT[911]      = 112'hC18F7320766F6C7574706174206D;
        inPKT[912]      = 112'hC190692073656420736167697474;
        inPKT[913]      = 112'hC19169732E0D0A0D0A4475697320;
        inPKT[914]      = 112'hC1926772617669646120656C656D;
        inPKT[915]      = 112'hC193656E74756D20696E74657264;
        inPKT[916]      = 112'hC194756D2E2050726F696E207369;
        inPKT[917]      = 112'hC1957420616D6574207175616D20;
        inPKT[918]      = 112'hC1966C6967756C612E2050686173;
        inPKT[919]      = 112'hC197656C6C757320636F6D6D6F64;
        inPKT[920]      = 112'hC1986F2C2075726E6120696E2063;
        inPKT[921]      = 112'hC1996F6E67756520766F6C757470;
        inPKT[922]      = 112'hC19A61742C206C6967756C612065;
        inPKT[923]      = 112'hC19B78207068617265747261206C;
        inPKT[924]      = 112'hC19C6967756C612C20696E206469;
        inPKT[925]      = 112'hC19D6374756D206D61676E61206F;
        inPKT[926]      = 112'hC19E726369206E6563206D617572;
        inPKT[927]      = 112'hC19F69732E204E756E6320617563;
        inPKT[928]      = 112'hC1A0746F7220636F6E7365637465;
        inPKT[929]      = 112'hC1A174757220766F6C7574706174;
        inPKT[930]      = 112'hC1A22E204D6F7262692074696E63;
        inPKT[931]      = 112'hC1A36964756E74206E6962682075;
        inPKT[932]      = 112'hC1A47420656E696D206566666963;
        inPKT[933]      = 112'hC1A5697475722067726176696461;
        inPKT[934]      = 112'hC1A62E2043757261626974757220;
        inPKT[935]      = 112'hC1A77669746165207175616D2065;
        inPKT[936]      = 112'hC1A8726F732E2044756973206672;
        inPKT[937]      = 112'hC1A9696E67696C6C612061632074;
        inPKT[938]      = 112'hC1AA6F72746F7220696E2074696E;
        inPKT[939]      = 112'hC1AB636964756E742E204E756E63;
        inPKT[940]      = 112'hC1AC2076656C206D617572697320;
        inPKT[941]      = 112'hC1AD72697375732E20446F6E6563;
        inPKT[942]      = 112'hC1AE20656C656966656E64206C69;
        inPKT[943]      = 112'hC1AF67756C612073616769747469;
        inPKT[944]      = 112'hC1B073206E6973692066696E6962;
        inPKT[945]      = 112'hC1B175732C2061207363656C6572;
        inPKT[946]      = 112'hC1B26973717565206C696265726F;
        inPKT[947]      = 112'hC1B32070656C6C656E7465737175;
        inPKT[948]      = 112'hC1B4652E20566573746962756C75;
        inPKT[949]      = 112'hC1B56D2074726973746971756520;
        inPKT[950]      = 112'hC1B66D61737361206E6962682C20;
        inPKT[951]      = 112'hC1B7617420766573746962756C75;
        inPKT[952]      = 112'hC1B86D206D61676E612066696E69;
        inPKT[953]      = 112'hC1B96275732065752E0D0A0D0A43;
        inPKT[954]      = 112'hC1BA757261626974757220696D70;
        inPKT[955]      = 112'hC1BB657264696574207075727573;
        inPKT[956]      = 112'hC1BC2065676574206E756E632075;
        inPKT[957]      = 112'hC1BD6C7472696365732C20766974;
        inPKT[958]      = 112'hC1BE61652076656E656E61746973;
        inPKT[959]      = 112'hC1BF206D6173736120636F6D6D6F;
        inPKT[960]      = 112'hC1C0646F2E2050656C6C656E7465;
        inPKT[961]      = 112'hC1C173717565206861626974616E;
        inPKT[962]      = 112'hC1C274206D6F7262692074726973;
        inPKT[963]      = 112'hC1C374697175652073656E656374;
        inPKT[964]      = 112'hC1C47573206574206E6574757320;
        inPKT[965]      = 112'hC1C56574206D616C657375616461;
        inPKT[966]      = 112'hC1C62066616D6573206163207475;
        inPKT[967]      = 112'hC1C7727069732065676573746173;
        inPKT[968]      = 112'hC1C82E20496E206665726D656E74;
        inPKT[969]      = 112'hC1C9756D2061742075726E61206E;
        inPKT[970]      = 112'hC1CA6F6E20636F6E76616C6C6973;
        inPKT[971]      = 112'hC1CB2E20446F6E65632061632061;
        inPKT[972]      = 112'hC1CC75677565206A7573746F2E20;
        inPKT[973]      = 112'hC1CD496E20617420656C69742065;
        inPKT[974]      = 112'hC1CE742061726375206D6178696D;
        inPKT[975]      = 112'hC1CF7573206C75637475732E2046;
        inPKT[976]      = 112'hC1D07573636520657569736D6F64;
        inPKT[977]      = 112'hC1D1206E756E63206E6563207665;
        inPKT[978]      = 112'hC1D26E656E617469732061756374;
        inPKT[979]      = 112'hC1D36F722E204C6F72656D206970;
        inPKT[980]      = 112'hC1D473756D20646F6C6F72207369;
        inPKT[981]      = 112'hC1D57420616D65742C20636F6E73;
        inPKT[982]      = 112'hC1D6656374657475722061646970;
        inPKT[983]      = 112'hC1D7697363696E6720656C69742E;
        inPKT[984]      = 112'hC1D820446F6E6563206469637475;
        inPKT[985]      = 112'hC1D96D2074656D706F7220727574;
        inPKT[986]      = 112'hC1DA72756D2E2053656420656C65;
        inPKT[987]      = 112'hC1DB6966656E64206469616D2069;
        inPKT[988]      = 112'hC1DC64206D6173736120696D7065;
        inPKT[989]      = 112'hC1DD72646965742C206163206F72;
        inPKT[990]      = 112'hC1DE6E617265206C696265726F20;
        inPKT[991]      = 112'hC1DF656C656966656E642E204D61;
        inPKT[992]      = 112'hC1E06563656E6173206F726E6172;
        inPKT[993]      = 112'hC1E165206D65747573206E756C6C;
        inPKT[994]      = 112'hC1E2612C2073697420616D657420;
        inPKT[995]      = 112'hC1E36665726D656E74756D20656C;
        inPKT[996]      = 112'hC1E4697420616C697175616D2069;
        inPKT[997]      = 112'hC1E5642E20446F6E656320756C74;
        inPKT[998]      = 112'hC1E6726963657320746F72746F72;
        inPKT[999]      = 112'hC1E720617420616E74652068656E;
        inPKT[1000]     = 112'hC1E86472657269742C2065752073;
        inPKT[1001]     = 112'hC1E961676974746973206A757374;
        inPKT[1002]     = 112'hC1EA6F20756C7472696365732E0D;
        inPKT[1003]     = 112'hC1EB0A0D0A5072616573656E7420;
        inPKT[1004]     = 112'hC1EC6C7563747573207072657469;
        inPKT[1005]     = 112'hC1ED756D206E657175652C207369;
        inPKT[1006]     = 112'hC1EE7420616D65742070656C6C65;
        inPKT[1007]     = 112'hC1EF6E746573717565206D617572;
        inPKT[1008]     = 112'hC1F0697320656C656D656E74756D;
        inPKT[1009]     = 112'hC1F1206E6F6E2E20557420626C61;
        inPKT[1010]     = 112'hC1F26E6469742070686172657472;
        inPKT[1011]     = 112'hC1F361206F64696F206E6F6E2065;
        inPKT[1012]     = 112'hC1F47569736D6F642E2051756973;
        inPKT[1013]     = 112'hC1F5717565207669746165206C65;
        inPKT[1014]     = 112'hC1F66F20616C697175616D2C2073;
        inPKT[1015]     = 112'hC1F76F64616C65732074656C6C75;
        inPKT[1016]     = 112'hC1F8732069642C20696163756C69;
        inPKT[1017]     = 112'hC1F973206D61757269732E204E61;
        inPKT[1018]     = 112'hC1FA6D2065666669636974757220;
        inPKT[1019]     = 112'hC1FB696E20707572757320736564;
        inPKT[1020]     = 112'hC1FC20616363756D73616E2E204D;
        inPKT[1021]     = 112'hC1FD616563656E61732073697420;
        inPKT[1022]     = 112'hC1FE616D65742063757273757320;
        inPKT[1023]     = 112'hC1FF66656C69732E205175697371;
        inPKT[1024]     = 112'hC10075652066617563696275732C;
        inPKT[1025]     = 112'hC101206475692065742061756374;
        inPKT[1026]     = 112'hC1026F72206C75637475732C2061;
        inPKT[1027]     = 112'hC1036E7465206572617420706F73;
        inPKT[1028]     = 112'hC104756572652065726F732C2075;
        inPKT[1029]     = 112'hC1057420636F6E76616C6C697320;
        inPKT[1030]     = 112'hC1066D65747573206C6563747573;
        inPKT[1031]     = 112'hC107207669746165206C656F2E20;
        inPKT[1032]     = 112'hC10853757370656E646973736520;
        inPKT[1033]     = 112'hC109706F74656E74692E20437261;
        inPKT[1034]     = 112'hC10A7320657420646F6C6F72206E;
        inPKT[1035]     = 112'hC10B6F6E2075726E61207363656C;
        inPKT[1036]     = 112'hC10C657269737175652074726973;
        inPKT[1037]     = 112'hC10D74697175652E204372617320;
        inPKT[1038]     = 112'hC10E72757472756D206E65632076;
        inPKT[1039]     = 112'hC10F656C69742061632073616769;
        inPKT[1040]     = 112'hC110747469732E20446F6E656320;
        inPKT[1041]     = 112'hC111656C656966656E642C206C61;
        inPKT[1042]     = 112'hC112637573207365642067726176;
        inPKT[1043]     = 112'hC113696461206D616C6573756164;
        inPKT[1044]     = 112'hC114612C20657820616E74652070;
        inPKT[1045]     = 112'hC1156C616365726174206C656374;
        inPKT[1046]     = 112'hC11675732C206567657420636F6E;
        inPKT[1047]     = 112'hC117677565206D61737361206D65;
        inPKT[1048]     = 112'hC118747573206964206C61637573;
        inPKT[1049]     = 112'hC1192E2053757370656E64697373;
        inPKT[1050]     = 112'hC11A652069642072757472756D20;
        inPKT[1051]     = 112'hC11B6C65637475732E2046757363;
        inPKT[1052]     = 112'hC11C65206D6178696D7573207365;
        inPKT[1053]     = 112'hC11D64206C6967756C6120736564;
        inPKT[1054]     = 112'hC11E20766976657272612E204E61;
        inPKT[1055]     = 112'hC11F6D206C756374757320646961;
        inPKT[1056]     = 112'hC1206D20616E74652C2076697461;
        inPKT[1057]     = 112'hC12165206F726E617265206E6571;
        inPKT[1058]     = 112'hC122756520766172697573206567;
        inPKT[1059]     = 112'hC12365742E0D0A0D0A50656C6C65;
        inPKT[1060]     = 112'hC1246E7465737175652061742065;
        inPKT[1061]     = 112'hC1256C6974206E6962682E205665;
        inPKT[1062]     = 112'hC12673746962756C756D20616E74;
        inPKT[1063]     = 112'hC1276520697073756D207072696D;
        inPKT[1064]     = 112'hC128697320696E20666175636962;
        inPKT[1065]     = 112'hC1297573206F726369206C756374;
        inPKT[1066]     = 112'hC12A757320657420756C74726963;
        inPKT[1067]     = 112'hC12B657320706F73756572652063;
        inPKT[1068]     = 112'hC12C7562696C6961204375726165;
        inPKT[1069]     = 112'hC12D3B2043757261626974757220;
        inPKT[1070]     = 112'hC12E666175636962757320646961;
        inPKT[1071]     = 112'hC12F6D206C656F2C206E65632065;
        inPKT[1072]     = 112'hC1307569736D6F642073656D2065;
        inPKT[1073]     = 112'hC13166666963697475722075742E;
        inPKT[1074]     = 112'hC132205574207665686963756C61;
        inPKT[1075]     = 112'hC133206175677565206163206C69;
        inPKT[1076]     = 112'hC1346265726F20696163756C6973;
        inPKT[1077]     = 112'hC1352C206E656320656C65696665;
        inPKT[1078]     = 112'hC1366E6420657820706F7274612E;
        inPKT[1079]     = 112'hC137204D6F7262692068656E6472;
        inPKT[1080]     = 112'hC138657269742067726176696461;
        inPKT[1081]     = 112'hC1392074696E636964756E742E20;
        inPKT[1082]     = 112'hC13A5072616573656E7420646F6C;
        inPKT[1083]     = 112'hC13B6F72206C616375732C207465;
        inPKT[1084]     = 112'hC13C6D707573206575206672696E;
        inPKT[1085]     = 112'hC13D67696C6C612073697420616D;
        inPKT[1086]     = 112'hC13E65742C20656C656966656E64;
        inPKT[1087]     = 112'hC13F20696E206E756C6C612E204E;
        inPKT[1088]     = 112'hC140756C6C61206D6F6C6C697320;
        inPKT[1089]     = 112'hC14165676574206D61676E61206E;
        inPKT[1090]     = 112'hC14265632068656E647265726974;
        inPKT[1091]     = 112'hC1432E20416C697175616D20636F;
        inPKT[1092]     = 112'hC1446E76616C6C69732073656D20;
        inPKT[1093]     = 112'hC14576697461652073617069656E;
        inPKT[1094]     = 112'hC1462064696374756D2C20757420;
        inPKT[1095]     = 112'hC147766573746962756C756D206C;
        inPKT[1096]     = 112'hC1486F72656D206672696E67696C;
        inPKT[1097]     = 112'hC1496C612E20446F6E6563207465;
        inPKT[1098]     = 112'hC14A6C6C7573206C696265726F2C;
        inPKT[1099]     = 112'hC14B206665756769617420757420;
        inPKT[1100]     = 112'hC14C66696E69627573206E65632C;
        inPKT[1101]     = 112'hC14D20616C697175616D20736974;
        inPKT[1102]     = 112'hC14E20616D6574206F7263692E20;
        inPKT[1103]     = 112'hC14F4E756E632073757363697069;
        inPKT[1104]     = 112'hC15074206E69736C206574206F72;
        inPKT[1105]     = 112'hC1516E6172652076657374696275;
        inPKT[1106]     = 112'hC1526C756D2E204E756C6C616D20;
        inPKT[1107]     = 112'hC1536C6F626F7274697320736170;
        inPKT[1108]     = 112'hC15469656E206A7573746F2C2073;
        inPKT[1109]     = 112'hC155697420616D6574206469676E;
        inPKT[1110]     = 112'hC156697373696D206E756C6C6120;
        inPKT[1111]     = 112'hC157636F6E64696D656E74756D20;
        inPKT[1112]     = 112'hC158696E2E20536564206D6F6C65;
        inPKT[1113]     = 112'hC1597374696520766F6C75747061;
        inPKT[1114]     = 112'hC15A74206E697369206174206665;
        inPKT[1115]     = 112'hC15B726D656E74756D2E204E756C;
        inPKT[1116]     = 112'hC15C6C61206D6F6C657374696520;
        inPKT[1117]     = 112'hC15D6E6973692073656420747572;
        inPKT[1118]     = 112'hC15E706973206D6F6C6573746965;
        inPKT[1119]     = 112'hC15F2C206E6F6E20696163756C69;
        inPKT[1120]     = 112'hC16073206E756E63206661756369;
        inPKT[1121]     = 112'hC1616275732E2041656E65616E20;
        inPKT[1122]     = 112'hC162696E74657264756D20706861;
        inPKT[1123]     = 112'hC163726574726120636F6E736563;
        inPKT[1124]     = 112'hC16474657475722E20457469616D;
        inPKT[1125]     = 112'hC165206578206F7263692C206961;
        inPKT[1126]     = 112'hC16663756C6973206E6F6E206575;
        inPKT[1127]     = 112'hC16769736D6F642069642C20756C;
        inPKT[1128]     = 112'hC1686C616D636F72706572207363;
        inPKT[1129]     = 112'hC169656C65726973717565206F64;
        inPKT[1130]     = 112'hC16A696F2E0D0A0D0A4E616D2075;
        inPKT[1131]     = 112'hC16B6C74726963657320656C6569;
        inPKT[1132]     = 112'hC16C66656E64206469616D2C2065;
        inPKT[1133]     = 112'hC16D67657420736F64616C657320;
        inPKT[1134]     = 112'hC16E73656D206D61747469732061;
        inPKT[1135]     = 112'hC16F632E2055742076656E656E61;
        inPKT[1136]     = 112'hC170746973206E69626820657520;
        inPKT[1137]     = 112'hC1716C65637475732074696E6369;
        inPKT[1138]     = 112'hC17264756E742064696374756D2E;
        inPKT[1139]     = 112'hC17320566976616D757320637572;
        inPKT[1140]     = 112'hC174737573206175677565207175;
        inPKT[1141]     = 112'hC1756973206C6F626F7274697320;
        inPKT[1142]     = 112'hC176657569736D6F642E204E756E;
        inPKT[1143]     = 112'hC1776320616C697175616D206469;
        inPKT[1144]     = 112'hC178616D20617420616E74652066;
        inPKT[1145]     = 112'hC1796163696C69736973206D6178;
        inPKT[1146]     = 112'hC17A696D75732E20457469616D20;
        inPKT[1147]     = 112'hC17B736564206C6F72656D206D61;
        inPKT[1148]     = 112'hC17C747469732C20636F6E76616C;
        inPKT[1149]     = 112'hC17D6C69732075726E6120766974;
        inPKT[1150]     = 112'hC17E61652C2074656D7075732073;
        inPKT[1151]     = 112'hC17F656D2E20566976616D757320;
        inPKT[1152]     = 112'hC1806567657374617320766F6C75;
        inPKT[1153]     = 112'hC181747061742065726F73206575;
        inPKT[1154]     = 112'hC18220756C7472696365732E2056;
        inPKT[1155]     = 112'hC1836573746962756C756D20756C;
        inPKT[1156]     = 112'hC1846C616D636F72706572206572;
        inPKT[1157]     = 112'hC1856174206E756E632C206E6F6E;
        inPKT[1158]     = 112'hC1862068656E647265726974206F;
        inPKT[1159]     = 112'hC18764696F2070656C6C656E7465;
        inPKT[1160]     = 112'hC188737175652069642E20467573;
        inPKT[1161]     = 112'hC18963652075726E612069707375;
        inPKT[1162]     = 112'hC18A6D2C206C6163696E69612069;
        inPKT[1163]     = 112'hC18B6E2073757363697069742076;
        inPKT[1164]     = 112'hC18C656C2C2073656D7065722069;
        inPKT[1165]     = 112'hC18D6E206F64696F2E2050656C6C;
        inPKT[1166]     = 112'hC18E656E74657371756520696420;
        inPKT[1167]     = 112'hC18F6E696268206E6973692E2041;
        inPKT[1168]     = 112'hC1906C697175616D20706F727461;
        inPKT[1169]     = 112'hC191206E69736C20657420657820;
        inPKT[1170]     = 112'hC192696163756C69732074726973;
        inPKT[1171]     = 112'hC19374697175652E20457469616D;
        inPKT[1172]     = 112'hC194206D61737361206F7263692C;
        inPKT[1173]     = 112'hC195206567657374617320736564;
        inPKT[1174]     = 112'hC196206C6F72656D20717569732C;
        inPKT[1175]     = 112'hC197206469676E697373696D2073;
        inPKT[1176]     = 112'hC198656D70657220616E74652E20;
        inPKT[1177]     = 112'hC19953757370656E646973736520;
        inPKT[1178]     = 112'hC19A74696E636964756E74206E69;
        inPKT[1179]     = 112'hC19B73692065782C207365642076;
        inPKT[1180]     = 112'hC19C6F6C75747061742065737420;
        inPKT[1181]     = 112'hC19D766172697573207669746165;
        inPKT[1182]     = 112'hC19E2E0D0A0D0A5365642073656D;
        inPKT[1183]     = 112'hC19F706572206C6163696E696120;
        inPKT[1184]     = 112'hC1A0646F6C6F722E204E616D2075;
        inPKT[1185]     = 112'hC1A1742076656C697420696E206C;
        inPKT[1186]     = 112'hC1A26163757320636F6E73656374;
        inPKT[1187]     = 112'hC1A36574757220636F6E76616C6C;
        inPKT[1188]     = 112'hC1A469732070656C6C656E746573;
        inPKT[1189]     = 112'hC1A5717565207365642073656D2E;
        inPKT[1190]     = 112'hC1A62053757370656E6469737365;
        inPKT[1191]     = 112'hC1A720636F6E64696D656E74756D;
        inPKT[1192]     = 112'hC1A820612065726F732069642075;
        inPKT[1193]     = 112'hC1A96C6C616D636F727065722E20;
        inPKT[1194]     = 112'hC1AA4D6F726269206C7563747573;
        inPKT[1195]     = 112'hC1AB2075726E612073697420616D;
        inPKT[1196]     = 112'hC1AC657420657569736D6F642069;
        inPKT[1197]     = 112'hC1AD6163756C69732E2050656C6C;
        inPKT[1198]     = 112'hC1AE656E74657371756520666163;
        inPKT[1199]     = 112'hC1AF696C69736973206D61757269;
        inPKT[1200]     = 112'hC1B07320657520656C656D656E74;
        inPKT[1201]     = 112'hC1B1756D207661726975732E204F;
        inPKT[1202]     = 112'hC1B272636920766172697573206E;
        inPKT[1203]     = 112'hC1B361746F7175652070656E6174;
        inPKT[1204]     = 112'hC1B469627573206574206D61676E;
        inPKT[1205]     = 112'hC1B5697320646973207061727475;
        inPKT[1206]     = 112'hC1B67269656E74206D6F6E746573;
        inPKT[1207]     = 112'hC1B72C206E617363657475722072;
        inPKT[1208]     = 112'hC1B869646963756C7573206D7573;
        inPKT[1209]     = 112'hC1B92E20446F6E6563206469676E;
        inPKT[1210]     = 112'hC1BA697373696D20612069707375;
        inPKT[1211]     = 112'hC1BB6D20756C7472696369657320;
        inPKT[1212]     = 112'hC1BC76656E656E617469732E2056;
        inPKT[1213]     = 112'hC1BD6976616D7573206E756E6320;
        inPKT[1214]     = 112'hC1BE76656C69742C207665686963;
        inPKT[1215]     = 112'hC1BF756C61207669746165206D61;
        inPKT[1216]     = 112'hC1C07373612075742C20636F6E76;
        inPKT[1217]     = 112'hC1C1616C6C697320636F6E736563;
        inPKT[1218]     = 112'hC1C2746574757220746F72746F72;
        inPKT[1219]     = 112'hC1C32E205175697371756520616C;
        inPKT[1220]     = 112'hC1C4697175616D2C206E69736C20;
        inPKT[1221]     = 112'hC1C5636F6E67756520626C616E64;
        inPKT[1222]     = 112'hC1C6697420756C74726963696573;
        inPKT[1223]     = 112'hC1C72C2075726E61207475727069;
        inPKT[1224]     = 112'hC1C873206D6174746973206D6167;
        inPKT[1225]     = 112'hC1C96E612C206E6F6E206665726D;
        inPKT[1226]     = 112'hC1CA656E74756D20647569207665;
        inPKT[1227]     = 112'hC1CB6C6974206575207175616D2E;
        inPKT[1228]     = 112'hC1CC0D0A0D0A496E207068617265;
        inPKT[1229]     = 112'hC1CD7472612076656C697420646F;
        inPKT[1230]     = 112'hC1CE6C6F722C2076697461652063;
        inPKT[1231]     = 112'hC1CF7572737573206F7263692066;
        inPKT[1232]     = 112'hC1D0696E696275732074696E6369;
        inPKT[1233]     = 112'hC1D164756E742E20566976616D75;
        inPKT[1234]     = 112'hC1D27320696420746F72746F7220;
        inPKT[1235]     = 112'hC1D372686F6E6375732C20736167;
        inPKT[1236]     = 112'hC1D46974746973206469616D2065;
        inPKT[1237]     = 112'hC1D56765742C207072657469756D;
        inPKT[1238]     = 112'hC1D6206D61757269732E20506861;
        inPKT[1239]     = 112'hC1D773656C6C757320656C656D65;
        inPKT[1240]     = 112'hC1D86E74756D20656E696D206665;
        inPKT[1241]     = 112'hC1D96C69732E204D617572697320;
        inPKT[1242]     = 112'hC1DA6575206E6571756520656765;
        inPKT[1243]     = 112'hC1DB742070757275732068656E64;
        inPKT[1244]     = 112'hC1DC726572697420677261766964;
        inPKT[1245]     = 112'hC1DD612E20416C697175616D206C;
        inPKT[1246]     = 112'hC1DE696265726F206E6962682C20;
        inPKT[1247]     = 112'hC1DF636F6E76616C6C6973206120;
        inPKT[1248]     = 112'hC1E06E69736C2065742C2068656E;
        inPKT[1249]     = 112'hC1E1647265726974207665737469;
        inPKT[1250]     = 112'hC1E262756C756D2066656C69732E;
        inPKT[1251]     = 112'hC1E320446F6E656320657569736D;
        inPKT[1252]     = 112'hC1E46F64206665726D656E74756D;
        inPKT[1253]     = 112'hC1E5207475727069732065752061;
        inPKT[1254]     = 112'hC1E67563746F722E2041656E6561;
        inPKT[1255]     = 112'hC1E76E20626962656E64756D2074;
        inPKT[1256]     = 112'hC1E8757270697320696E206F6469;
        inPKT[1257]     = 112'hC1E96F20636F6E76616C6C69732C;
        inPKT[1258]     = 112'hC1EA207669746165207661726975;
        inPKT[1259]     = 112'hC1EB73206578206C616F72656574;
        inPKT[1260]     = 112'hC1EC2E2046757363652076656C20;
        inPKT[1261]     = 112'hC1ED6D6920766974616520646F6C;
        inPKT[1262]     = 112'hC1EE6F7220666575676961742076;
        inPKT[1263]     = 112'hC1EF756C707574617465206E6563;
        inPKT[1264]     = 112'hC1F0207574206E756E632E204372;
        inPKT[1265]     = 112'hC1F1617320646170696275732C20;
        inPKT[1266]     = 112'hC1F2616E74652069642076656869;
        inPKT[1267]     = 112'hC1F363756C6120616C697175616D;
        inPKT[1268]     = 112'hC1F42C20656C69742065726F7320;
        inPKT[1269]     = 112'hC1F57361676974746973206D692C;
        inPKT[1270]     = 112'hC1F6206E6F6E20656C656966656E;
        inPKT[1271]     = 112'hC1F764206578206E756C6C612065;
        inPKT[1272]     = 112'hC1F86765742076656C69742E2053;
        inPKT[1273]     = 112'hC1F9757370656E64697373652069;
        inPKT[1274]     = 112'hC1FA64206469616D206475692E20;
        inPKT[1275]     = 112'hC1FB53757370656E646973736520;
        inPKT[1276]     = 112'hC1FC7072657469756D206A757374;
        inPKT[1277]     = 112'hC1FD6F20736564206E6962682070;
        inPKT[1278]     = 112'hC1FE6F72747469746F722C207665;
        inPKT[1279]     = 112'hC1FF6C20696E74657264756D206D;
        inPKT[1280]     = 112'hC1006175726973206D6178696D75;
        inPKT[1281]     = 112'hC101732E20557420616C69717561;
        inPKT[1282]     = 112'hC1026D206C616375732070757275;
        inPKT[1283]     = 112'hC103732C2073697420616D657420;
        inPKT[1284]     = 112'hC104696D70657264696574206E69;
        inPKT[1285]     = 112'hC105626820666575676961742069;
        inPKT[1286]     = 112'hC106642E20496E7465676572206C;
        inPKT[1287]     = 112'hC1076F72656D206D61757269732C;
        inPKT[1288]     = 112'hC108207072657469756D206E6F6E;
        inPKT[1289]     = 112'hC109206E6973692065742C206461;
        inPKT[1290]     = 112'hC10A70696275732066696E696275;
        inPKT[1291]     = 112'hC10B73206F7263692E0D0A0D0A56;
        inPKT[1292]     = 112'hC10C6573746962756C756D206961;
        inPKT[1293]     = 112'hC10D63756C69732C206D61676E61;
        inPKT[1294]     = 112'hC10E206174206D6174746973206D;
        inPKT[1295]     = 112'hC10F6178696D75732C2061726375;
        inPKT[1296]     = 112'hC110206572617420646170696275;
        inPKT[1297]     = 112'hC11173206E756E632C2061207661;
        inPKT[1298]     = 112'hC11272697573206D657475732066;
        inPKT[1299]     = 112'hC113656C697320736564206F7263;
        inPKT[1300]     = 112'hC114692E204E756C6C616D206D69;
        inPKT[1301]     = 112'hC115206E6962682C20656C656966;
        inPKT[1302]     = 112'hC116656E64206E656320756C7472;
        inPKT[1303]     = 112'hC11769636573206E65632C20636F;
        inPKT[1304]     = 112'hC1186E7365637465747572206163;
        inPKT[1305]     = 112'hC11920656E696D2E20536564206C;
        inPKT[1306]     = 112'hC11A75637475732073656D207175;
        inPKT[1307]     = 112'hC11B69732074656D706F7220636F;
        inPKT[1308]     = 112'hC11C6E6775652E2053757370656E;
        inPKT[1309]     = 112'hC11D646973736520706F74656E74;
        inPKT[1310]     = 112'hC11E692E20457469616D20656765;
        inPKT[1311]     = 112'hC11F74206C696265726F2076656C;
        inPKT[1312]     = 112'hC12069742E204475697320766573;
        inPKT[1313]     = 112'hC121746962756C756D20636F6E73;
        inPKT[1314]     = 112'hC122657175617420706F7274612E;
        inPKT[1315]     = 112'hC123204D617572697320706F7274;
        inPKT[1316]     = 112'hC1247469746F7220747572706973;
        inPKT[1317]     = 112'hC12520696E206D6173736120616C;
        inPKT[1318]     = 112'hC126697175616D20636F6E677565;
        inPKT[1319]     = 112'hC1272E204E756C6C6120636F6E73;
        inPKT[1320]     = 112'hC128656374657475722075726E61;
        inPKT[1321]     = 112'hC129206D657475732C2069642069;
        inPKT[1322]     = 112'hC12A6163756C6973206E756E6320;
        inPKT[1323]     = 112'hC12B756C74726963696573206567;
        inPKT[1324]     = 112'hC12C65742E204375726162697475;
        inPKT[1325]     = 112'hC12D72206D6175726973206E6571;
        inPKT[1326]     = 112'hC12E75652C20626962656E64756D;
        inPKT[1327]     = 112'hC12F207365642065726F73206174;
        inPKT[1328]     = 112'hC1302C206D6178696D757320756C;
        inPKT[1329]     = 112'hC131747269636573207475727069;
        inPKT[1330]     = 112'hC132732E0D0A496E74657264756D;
        inPKT[1331]     = 112'hC133206574206D616C6573756164;
        inPKT[1332]     = 112'hC134612066616D65732061632061;
        inPKT[1333]     = 112'hC1356E746520697073756D207072;
        inPKT[1334]     = 112'hC136696D697320696E2066617563;
        inPKT[1335]     = 112'hC137696275732E2050656C6C656E;
        inPKT[1336]     = 112'hC13874657371756520736F6C6C69;
        inPKT[1337]     = 112'hC1396369747564696E20626C616E;
        inPKT[1338]     = 112'hC13A646974206665726D656E7475;
        inPKT[1339]     = 112'hC13B6D2E2050656C6C656E746573;
        inPKT[1340]     = 112'hC13C717565206E6F6E206C696775;
        inPKT[1341]     = 112'hC13D6C6120657520657261742076;
        inPKT[1342]     = 112'hC13E656E656E6174697320657569;
        inPKT[1343]     = 112'hC13F736D6F642E2050656C6C656E;
        inPKT[1344]     = 112'hC14074657371756520736F64616C;
        inPKT[1345]     = 112'hC141657320766573746962756C75;
        inPKT[1346]     = 112'hC1426D20636F6E76616C6C69732E;
        inPKT[1347]     = 112'hC1432050726F696E206D6F6C6573;
        inPKT[1348]     = 112'hC144746965207072657469756D20;
        inPKT[1349]     = 112'hC14565726F732076656C20656765;
        inPKT[1350]     = 112'hC146737461732E204D6F72626920;
        inPKT[1351]     = 112'hC147736F6C6C696369747564696E;
        inPKT[1352]     = 112'hC148207075727573206163206665;
        inPKT[1353]     = 112'hC149726D656E74756D206D617474;
        inPKT[1354]     = 112'hC14A69732E204E756E632076656C;
        inPKT[1355]     = 112'hC14B2074696E636964756E74206C;
        inPKT[1356]     = 112'hC14C696265726F2E204E756C6C61;
        inPKT[1357]     = 112'hC14D20616C697175657420697073;
        inPKT[1358]     = 112'hC14E756D206E6563207175616D20;
        inPKT[1359]     = 112'hC14F696D7065726469657420696E;
        inPKT[1360]     = 112'hC15074657264756D2E2050726165;
        inPKT[1361]     = 112'hC15173656E74206C6967756C6120;
        inPKT[1362]     = 112'hC15266656C69732C20696163756C;
        inPKT[1363]     = 112'hC153697320617420616C69717565;
        inPKT[1364]     = 112'hC154742061742C20736167697474;
        inPKT[1365]     = 112'hC1556973207175697320656C6974;
        inPKT[1366]     = 112'hC1562E0D0A517569737175652076;
        inPKT[1367]     = 112'hC157656C20696D70657264696574;
        inPKT[1368]     = 112'hC158206E6962682E205068617365;
        inPKT[1369]     = 112'hC1596C6C75732072757472756D20;
        inPKT[1370]     = 112'hC15A6469676E697373696D207269;
        inPKT[1371]     = 112'hC15B737573206E6F6E2074696E63;
        inPKT[1372]     = 112'hC15C6964756E742E205665737469;
        inPKT[1373]     = 112'hC15D62756C756D206E756E632069;
        inPKT[1374]     = 112'hC15E7073756D2C2076656E656E61;
        inPKT[1375]     = 112'hC15F746973206567657420706F72;
        inPKT[1376]     = 112'hC160746120696E2C20636F6E7365;
        inPKT[1377]     = 112'hC161637465747572206575206572;
        inPKT[1378]     = 112'hC16261742E20446F6E6563207665;
        inPKT[1379]     = 112'hC163686963756C6120616E746520;
        inPKT[1380]     = 112'hC16476656C2072686F6E63757320;
        inPKT[1381]     = 112'hC16566617563696275732E205065;
        inPKT[1382]     = 112'hC1666C6C656E746573717565206A;
        inPKT[1383]     = 112'hC1677573746F20746F72746F722C;
        inPKT[1384]     = 112'hC16820766F6C757470617420696E;
        inPKT[1385]     = 112'hC169206D61757269732061742C20;
        inPKT[1386]     = 112'hC16A766172697573207068617265;
        inPKT[1387]     = 112'hC16B7472612072697375732E2051;
        inPKT[1388]     = 112'hC16C756973717565207574206469;
        inPKT[1389]     = 112'hC16D616D2073757363697069742C;
        inPKT[1390]     = 112'hC16E20736F6C6C69636974756469;
        inPKT[1391]     = 112'hC16F6E2073617069656E2065742C;
        inPKT[1392]     = 112'hC17020696E74657264756D206C61;
        inPKT[1393]     = 112'hC1716375732E204D6F7262692072;
        inPKT[1394]     = 112'hC172697375732073656D2C207065;
        inPKT[1395]     = 112'hC1736C6C656E7465737175652065;
        inPKT[1396]     = 112'hC174742074757270697320696E2C;
        inPKT[1397]     = 112'hC17520626C616E64697420736F6C;
        inPKT[1398]     = 112'hC1766C696369747564696E207365;
        inPKT[1399]     = 112'hC1776D2E20536564206566666963;
        inPKT[1400]     = 112'hC17869747572206C696265726F20;
        inPKT[1401]     = 112'hC17971756973207072657469756D;
        inPKT[1402]     = 112'hC17A207072657469756D2E204E75;
        inPKT[1403]     = 112'hC17B6C6C616D20617563746F7220;
        inPKT[1404]     = 112'hC17C7361676974746973206C6F72;
        inPKT[1405]     = 112'hC17D656D2C20616320756C747269;
        inPKT[1406]     = 112'hC17E6365732061726375206D6178;
        inPKT[1407]     = 112'hC17F696D757320656765742E0D0A;
        inPKT[1408]     = 112'hC180566573746962756C756D2076;
        inPKT[1409]     = 112'hC1816F6C7574706174206C696775;
        inPKT[1410]     = 112'hC1826C6120617563746F72207365;
        inPKT[1411]     = 112'hC1836D20766976657272612C2075;
        inPKT[1412]     = 112'hC1846C6C616D636F727065722065;
        inPKT[1413]     = 112'hC1857569736D6F64206E65717565;
        inPKT[1414]     = 112'hC18620706F72747469746F722E20;
        inPKT[1415]     = 112'hC18753757370656E646973736520;
        inPKT[1416]     = 112'hC18876697665727261207363656C;
        inPKT[1417]     = 112'hC18965726973717565206F64696F;
        inPKT[1418]     = 112'hC18A2072686F6E63757320766F6C;
        inPKT[1419]     = 112'hC18B75747061742E20416C697175;
        inPKT[1420]     = 112'hC18C616D206572617420766F6C75;
        inPKT[1421]     = 112'hC18D747061742E2053757370656E;
        inPKT[1422]     = 112'hC18E646973736520706F74656E74;
        inPKT[1423]     = 112'hC18F692E20496E20686163206861;
        inPKT[1424]     = 112'hC1906269746173736520706C6174;
        inPKT[1425]     = 112'hC19165612064696374756D73742E;
        inPKT[1426]     = 112'hC1922050726F696E207574206E75;
        inPKT[1427]     = 112'hC1936C6C61207574206475692073;
        inPKT[1428]     = 112'hC19463656C657269737175652064;
        inPKT[1429]     = 112'hC195696374756D2E205175697371;
        inPKT[1430]     = 112'hC196756520737573636970697420;
        inPKT[1431]     = 112'hC1976E69626820706F7375657265;
        inPKT[1432]     = 112'hC198207175616D2076756C707574;
        inPKT[1433]     = 112'hC1996174652C206575206C616369;
        inPKT[1434]     = 112'hC19A6E696120616E746520677261;
        inPKT[1435]     = 112'hC19B766964612E20437572616269;
        inPKT[1436]     = 112'hC19C747572206D61737361206C6F;
        inPKT[1437]     = 112'hC19D72656D2C206F726E61726520;
        inPKT[1438]     = 112'hC19E6575206D6F6C6C6973206174;
        inPKT[1439]     = 112'hC19F2C207068617265747261206E;
        inPKT[1440]     = 112'hC1A06563206D617373612E204E75;
        inPKT[1441]     = 112'hC1A16C6C612066696E6962757320;
        inPKT[1442]     = 112'hC1A2656C656966656E64206F7263;
        inPKT[1443]     = 112'hC1A3692073697420616D65742063;
        inPKT[1444]     = 112'hC1A46F6E73656374657475722E20;
        inPKT[1445]     = 112'hC1A55365642074656D7075732076;
        inPKT[1446]     = 112'hC1A6697461652061726375206E65;
        inPKT[1447]     = 112'hC1A763206665726D656E74756D2E;
        inPKT[1448]     = 112'hC1A82041656E65616E2070656C6C;
        inPKT[1449]     = 112'hC1A9656E74657371756520766974;
        inPKT[1450]     = 112'hC1AA616520646F6C6F7220696E20;
        inPKT[1451]     = 112'hC1AB616363756D73616E2E204372;
        inPKT[1452]     = 112'hC1AC6173206469676E697373696D;
        inPKT[1453]     = 112'hC1AD2076756C707574617465206D;
        inPKT[1454]     = 112'hC1AE6F6C6C69732E204D61757269;
        inPKT[1455]     = 112'hC1AF7320706F7274612076656E65;
        inPKT[1456]     = 112'hC1B06E617469732072697375732C;
        inPKT[1457]     = 112'hC1B1206575207472697374697175;
        inPKT[1458]     = 112'hC1B26520646F6C6F722072757472;
        inPKT[1459]     = 112'hC1B3756D20696E2E204675736365;
        inPKT[1460]     = 112'hC1B420636F6E64696D656E74756D;
        inPKT[1461]     = 112'hC1B5206F7263692066656C69732C;
        inPKT[1462]     = 112'hC1B62073697420616D657420636F;
        inPKT[1463]     = 112'hC1B76E76616C6C6973206C696265;
        inPKT[1464]     = 112'hC1B8726F2074696E636964756E74;
        inPKT[1465]     = 112'hC1B92061632E0D0A566573746962;
        inPKT[1466]     = 112'hC1BA756C756D20696D7065726469;
        inPKT[1467]     = 112'hC1BB657420656C69742074656D70;
        inPKT[1468]     = 112'hC1BC6F72207175616D2067726176;
        inPKT[1469]     = 112'hC1BD6964612C207574206D616C65;
        inPKT[1470]     = 112'hC1BE73756164612074656C6C7573;
        inPKT[1471]     = 112'hC1BF20696D706572646965742E20;
        inPKT[1472]     = 112'hC1C050686173656C6C7573206F64;
        inPKT[1473]     = 112'hC1C1696F2073656D2C206D617474;
        inPKT[1474]     = 112'hC1C269732073656420756C747269;
        inPKT[1475]     = 112'hC1C36365732061742C2076697665;
        inPKT[1476]     = 112'hC1C47272612076656C206475692E;
        inPKT[1477]     = 112'hC1C5204E756E632075726E61206D;
        inPKT[1478]     = 112'hC1C6657475732C206C7563747573;
        inPKT[1479]     = 112'hC1C7206163206D6178696D757320;
        inPKT[1480]     = 112'hC1C8696E2C20636F6E7365637465;
        inPKT[1481]     = 112'hC1C9747572206E6F6E206E697369;
        inPKT[1482]     = 112'hC1CA2E204E756C6C612073697420;
        inPKT[1483]     = 112'hC1CB616D657420626962656E6475;
        inPKT[1484]     = 112'hC1CC6D2076656C69742E20446F6E;
        inPKT[1485]     = 112'hC1CD6563207175697320656E696D;
        inPKT[1486]     = 112'hC1CE206E6F6E2072697375732062;
        inPKT[1487]     = 112'hC1CF6C616E64697420666163696C;
        inPKT[1488]     = 112'hC1D0697369732071756973206E65;
        inPKT[1489]     = 112'hC1D1632072697375732E20437572;
        inPKT[1490]     = 112'hC1D2616269747572206575206573;
        inPKT[1491]     = 112'hC1D374207669746165206C656374;
        inPKT[1492]     = 112'hC1D4757320626C616E6469742061;
        inPKT[1493]     = 112'hC1D56C69717565742E2056657374;
        inPKT[1494]     = 112'hC1D66962756C756D20616E746520;
        inPKT[1495]     = 112'hC1D7697073756D207072696D6973;
        inPKT[1496]     = 112'hC1D820696E206661756369627573;
        inPKT[1497]     = 112'hC1D9206F726369206C7563747573;
        inPKT[1498]     = 112'hC1DA20657420756C747269636573;
        inPKT[1499]     = 112'hC1DB20706F737565726520637562;
        inPKT[1500]     = 112'hC1DC696C69612043757261653B20;
        inPKT[1501]     = 112'hC1DD566573746962756C756D2061;
        inPKT[1502]     = 112'hC1DE63206469676E697373696D20;
        inPKT[1503]     = 112'hC1DF6E756E632E20517569737175;
        inPKT[1504]     = 112'hC1E06520696E2073616769747469;
        inPKT[1505]     = 112'hC1E1732074656C6C75732C207369;
        inPKT[1506]     = 112'hC1E27420616D6574206665726D65;
        inPKT[1507]     = 112'hC1E36E74756D206E6962682E0D0A;
        inPKT[1508]     = 112'hC1E4496E206469676E697373696D;
        inPKT[1509]     = 112'hC1E5207269737573207669746165;
        inPKT[1510]     = 112'hC1E6207075727573207665737469;
        inPKT[1511]     = 112'hC1E762756C756D2C20617420656C;
        inPKT[1512]     = 112'hC1E8656D656E74756D206E756C6C;
        inPKT[1513]     = 112'hC1E96120706F73756572652E2053;
        inPKT[1514]     = 112'hC1EA6564206D6174746973206E75;
        inPKT[1515]     = 112'hC1EB6E63206E6962682E20537573;
        inPKT[1516]     = 112'hC1EC70656E64697373652070656C;
        inPKT[1517]     = 112'hC1ED6C656E74657371756520706C;
        inPKT[1518]     = 112'hC1EE616365726174207363656C65;
        inPKT[1519]     = 112'hC1EF7269737175652E2041656E65;
        inPKT[1520]     = 112'hC1F0616E2066657567696174206D;
        inPKT[1521]     = 112'hC1F1617572697320696420636F6E;
        inPKT[1522]     = 112'hC1F2677565206C6163696E69612E;
        inPKT[1523]     = 112'hC1F320457469616D207375736369;
        inPKT[1524]     = 112'hC1F4706974206C6967756C612074;
        inPKT[1525]     = 112'hC1F5656C6C75732C206120636F6E;
        inPKT[1526]     = 112'hC1F6677565206C65637475732061;
        inPKT[1527]     = 112'hC1F76C697175616D207665686963;
        inPKT[1528]     = 112'hC1F8756C612E2053757370656E64;
        inPKT[1529]     = 112'hC1F969737365206567657420616E;
        inPKT[1530]     = 112'hC1FA74652076656C20656E696D20;
        inPKT[1531]     = 112'hC1FB6D616C657375616461207669;
        inPKT[1532]     = 112'hC1FC76657272612E2050726F696E;
        inPKT[1533]     = 112'hC1FD2074696E636964756E742061;
        inPKT[1534]     = 112'hC1FE72637520656765742076756C;
        inPKT[1535]     = 112'hC1FF70757461746520616363756D;
        inPKT[1536]     = 112'hC10073616E2E20496E2076697461;
        inPKT[1537]     = 112'hC10165206469616D206E6962682E;
        inPKT[1538]     = 112'hC102204D6F726269206D6178696D;
        inPKT[1539]     = 112'hC10375732066656C697320696420;
        inPKT[1540]     = 112'hC104636F6E736563746574757220;
        inPKT[1541]     = 112'hC105616C697175616D2E204E756C;
        inPKT[1542]     = 112'hC1066C6120666163696C6973692E;
        inPKT[1543]     = 112'hC1070D0A566573746962756C756D;
        inPKT[1544]     = 112'hC10820766573746962756C756D20;
        inPKT[1545]     = 112'hC10965666669636974757220746F;
        inPKT[1546]     = 112'hC10A72746F722073697420616D65;
        inPKT[1547]     = 112'hC10B7420666163696C697369732E;
        inPKT[1548]     = 112'hC10C204D616563656E6173206E6F;
        inPKT[1549]     = 112'hC10D6E2074656C6C7573206F7263;
        inPKT[1550]     = 112'hC10E692E2050686173656C6C7573;
        inPKT[1551]     = 112'hC10F206E6F6E206C756374757320;
        inPKT[1552]     = 112'hC1106A7573746F2C206174207375;
        inPKT[1553]     = 112'hC1117363697069742074656C6C75;
        inPKT[1554]     = 112'hC112732E2046757363652068656E;
        inPKT[1555]     = 112'hC113647265726974206E6563206E;
        inPKT[1556]     = 112'hC1146962682076656C2063757273;
        inPKT[1557]     = 112'hC11575732E2053757370656E6469;
        inPKT[1558]     = 112'hC11673736520706F74656E74692E;
        inPKT[1559]     = 112'hC1172044756973206C6967756C61;
        inPKT[1560]     = 112'hC1182066656C69732C2065666669;
        inPKT[1561]     = 112'hC11963697475722065742076656C;
        inPKT[1562]     = 112'hC11A69742061742C20666163696C;
        inPKT[1563]     = 112'hC11B6973697320636F6E76616C6C;
        inPKT[1564]     = 112'hC11C6973206A7573746F2E204E75;
        inPKT[1565]     = 112'hC11D6C6C616D206C6F626F727469;
        inPKT[1566]     = 112'hC11E732070656C6C656E74657371;
        inPKT[1567]     = 112'hC11F756520736F6C6C6963697475;
        inPKT[1568]     = 112'hC12064696E2E204E616D20736974;
        inPKT[1569]     = 112'hC12120616D657420646F6C6F7220;
        inPKT[1570]     = 112'hC12273697420616D6574206C6563;
        inPKT[1571]     = 112'hC12374757320696D706572646965;
        inPKT[1572]     = 112'hC1247420636F6E7365717561742E;
        inPKT[1573]     = 112'hC12520416C697175616D206C7563;
        inPKT[1574]     = 112'hC126747573207363656C65726973;
        inPKT[1575]     = 112'hC1277175652070757275732C2069;
        inPKT[1576]     = 112'hC12864206672696E67696C6C6120;
        inPKT[1577]     = 112'hC12973656D20766F6C7574706174;
        inPKT[1578]     = 112'hC12A2061632E205365642074656D;
        inPKT[1579]     = 112'hC12B706F722C20656E696D206567;
        inPKT[1580]     = 112'hC12C657420657569736D6F642066;
        inPKT[1581]     = 112'hC12D6163696C697369732C206E69;
        inPKT[1582]     = 112'hC12E73692065782073656D706572;
        inPKT[1583]     = 112'hC12F20697073756D2C20696E2073;
        inPKT[1584]     = 112'hC13061676974746973206F726369;
        inPKT[1585]     = 112'hC131207175616D20696E206C6563;
        inPKT[1586]     = 112'hC1327475732E2055742076697461;
        inPKT[1587]     = 112'hC1336520656C6974206C6967756C;
        inPKT[1588]     = 112'hC134612E204E756E632065676573;
        inPKT[1589]     = 112'hC1357461732C206D692076697461;
        inPKT[1590]     = 112'hC1366520696163756C6973206D61;
        inPKT[1591]     = 112'hC137747469732C20647569206E69;
        inPKT[1592]     = 112'hC138626820656C656966656E6420;
        inPKT[1593]     = 112'hC1396E69736C2C20656765742070;
        inPKT[1594]     = 112'hC13A6F727461206C696265726F20;
        inPKT[1595]     = 112'hC13B617567756520717569732065;
        inPKT[1596]     = 112'hC13C6E696D2E2053656420736974;
        inPKT[1597]     = 112'hC13D20616D65742070756C76696E;
        inPKT[1598]     = 112'hC13E61722065782C2076656C2070;
        inPKT[1599]     = 112'hC13F656C6C656E74657371756520;
        inPKT[1600]     = 112'hC1406C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
