`include "SIMON_defintions.svh"

module test_SIMON_9696_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 800
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 208'hE5000D0C0B0A0908050403020100000000000000000000000000;
        inPKT[1]        = 208'hC5014C6F72656D20697073756D20646F6C6F722073697420616D;
        inPKT[2]        = 208'hC50265742C20636F6E7365637465747572206164697069736369;
        inPKT[3]        = 208'hC5036E6720656C69742E2043757261626974757220756C6C616D;
        inPKT[4]        = 208'hC504636F727065722074656D707573206E6973692C2065742070;
        inPKT[5]        = 208'hC5056F73756572652075726E612E2041656E65616E2073656420;
        inPKT[6]        = 208'hC50667726176696461206C616375732E204E756C6C6120666163;
        inPKT[7]        = 208'hC507696C6973692E204E756C6C612074656D707573206F726369;
        inPKT[8]        = 208'hC508207175697320656C697420666575676961742C2076656C20;
        inPKT[9]        = 208'hC50973656D706572206C656F20696D706572646965742E204D61;
        inPKT[10]       = 208'hC50A6563656E6173206574206E756E6320696E206E6962682066;
        inPKT[11]       = 208'hC50B6163696C6973697320636F6E76616C6C69732E2053656420;
        inPKT[12]       = 208'hC50C636F6E6775652068656E64726572697420696163756C6973;
        inPKT[13]       = 208'hC50D2E20566976616D7573207665686963756C61206C75637475;
        inPKT[14]       = 208'hC50E73206573742C207669746165207375736369706974206E69;
        inPKT[15]       = 208'hC50F736C20706F72747469746F722061632E0D0A0D0A446F6E65;
        inPKT[16]       = 208'hC51063206D6F6C65737469652073617069656E2069642076756C;
        inPKT[17]       = 208'hC51170757461746520766573746962756C756D2E204E756C6C61;
        inPKT[18]       = 208'hC51220696E206C6967756C61206672696E67696C6C612C20756C;
        inPKT[19]       = 208'hC5136C616D636F727065722075726E612065742C20706F727474;
        inPKT[20]       = 208'hC51469746F72206C65637475732E205175697371756520626C61;
        inPKT[21]       = 208'hC5156E646974206575206D61757269732061632068656E647265;
        inPKT[22]       = 208'hC5167269742E204E756C6C612076656E656E617469732C206D65;
        inPKT[23]       = 208'hC517747573206574206C7563747573206672696E67696C6C612C;
        inPKT[24]       = 208'hC518206E6962682076656C697420756C6C616D636F7270657220;
        inPKT[25]       = 208'hC5196469616D2C20656765742065666669636974757220697073;
        inPKT[26]       = 208'hC51A756D20747572706973206174206E6962682E205574206567;
        inPKT[27]       = 208'hC51B6574207072657469756D2065726F732C2065676574206469;
        inPKT[28]       = 208'hC51C6374756D206C616375732E204D616563656E617320757420;
        inPKT[29]       = 208'hC51D656E696D2065782E2041656E65616E207669746165207365;
        inPKT[30]       = 208'hC51E6D7065722066656C69732C2073656420756C747269636965;
        inPKT[31]       = 208'hC51F732072697375732E20446F6E656320636F6E736563746574;
        inPKT[32]       = 208'hC5207572206D69206E69736C2C20617420637572737573206970;
        inPKT[33]       = 208'hC52173756D206772617669646120612E2050686173656C6C7573;
        inPKT[34]       = 208'hC5222073697420616D6574206D61676E612076656C2069707375;
        inPKT[35]       = 208'hC5236D206567657374617320706F7274612E20566976616D7573;
        inPKT[36]       = 208'hC524206C756374757320656E696D20656765742074656D706F72;
        inPKT[37]       = 208'hC5252073616769747469732E20416C697175616D20626962656E;
        inPKT[38]       = 208'hC52664756D2073656D206120636F6E7365637465747572206566;
        inPKT[39]       = 208'hC527666963697475722E20446F6E6563207363656C6572697371;
        inPKT[40]       = 208'hC528756520616C697175616D206375727375732E204375726162;
        inPKT[41]       = 208'hC529697475722073697420616D657420626962656E64756D2065;
        inPKT[42]       = 208'hC52A6C69742E20536564206469616D206A7573746F2C20696163;
        inPKT[43]       = 208'hC52B756C69732071756973206E756C6C612076697461652C2061;
        inPKT[44]       = 208'hC52C6C697175616D20657569736D6F642066656C69732E0D0A0D;
        inPKT[45]       = 208'hC52D0A50726F696E20646170696275732C206469616D2076756C;
        inPKT[46]       = 208'hC52E707574617465206672696E67696C6C61206D616C65737561;
        inPKT[47]       = 208'hC52F64612C206A7573746F20707572757320636F6D6D6F646F20;
        inPKT[48]       = 208'hC530646F6C6F722C2075742064696374756D2065726174206E75;
        inPKT[49]       = 208'hC5316E632072757472756D2075726E612E204E756C6C61206772;
        inPKT[50]       = 208'hC53261766964612075726E6120766974616520696D7065726469;
        inPKT[51]       = 208'hC5336574206C616F726565742E2050656C6C656E746573717565;
        inPKT[52]       = 208'hC5342072686F6E63757320626962656E64756D206E6962682C20;
        inPKT[53]       = 208'hC5356964206D6F6C6C6973206469616D20737573636970697420;
        inPKT[54]       = 208'hC53661632E2050656C6C656E7465737175652076656C20696163;
        inPKT[55]       = 208'hC537756C6973206475692E204D6F72626920617420616C697175;
        inPKT[56]       = 208'hC5386574206D617373612E2050726F696E207669746165206F72;
        inPKT[57]       = 208'hC5396E617265206F64696F2C2065752076756C70757461746520;
        inPKT[58]       = 208'hC53A697073756D2E2050726F696E206C6F626F727469732C2073;
        inPKT[59]       = 208'hC53B656D206E656320657569736D6F642074696E636964756E74;
        inPKT[60]       = 208'hC53C2C206175677565206D6175726973207363656C6572697371;
        inPKT[61]       = 208'hC53D7565206D61676E612C20657420706F7375657265206D6920;
        inPKT[62]       = 208'hC53E6E69736C206E6563206E6973692E20467573636520656C69;
        inPKT[63]       = 208'hC53F74206E657175652C20766172697573206574206672696E67;
        inPKT[64]       = 208'hC540696C6C612076697461652C207661726975732076656C206E;
        inPKT[65]       = 208'hC541657175652E204E756C6C612065742074656D707573206A75;
        inPKT[66]       = 208'hC54273746F2E204D6F72626920756C6C616D636F727065722073;
        inPKT[67]       = 208'hC5437573636970697420636F6E6775652E2053656420656C6569;
        inPKT[68]       = 208'hC54466656E64206F64696F206163207375736369706974206469;
        inPKT[69]       = 208'hC545676E697373696D2E205175697371756520616E746520656E;
        inPKT[70]       = 208'hC546696D2C20626C616E64697420696E20636F6E736571756174;
        inPKT[71]       = 208'hC5472061632C20696E74657264756D2076697461652070757275;
        inPKT[72]       = 208'hC548732E204D617572697320657569736D6F6420706F73756572;
        inPKT[73]       = 208'hC54965206C65637475732E20566976616D757320696E74657264;
        inPKT[74]       = 208'hC54A756D207175616D2065752073656D70657220666175636962;
        inPKT[75]       = 208'hC54B75732E0D0A0D0A496E206D6F6C6573746965206E756C6C61;
        inPKT[76]       = 208'hC54C20616E74652C20616320696E74657264756D206D61676E61;
        inPKT[77]       = 208'hC54D20636F6E64696D656E74756D20636F6E64696D656E74756D;
        inPKT[78]       = 208'hC54E2E204475697320756C7472696369657320736F64616C6573;
        inPKT[79]       = 208'hC54F206E756C6C612C2073697420616D657420756C6C616D636F;
        inPKT[80]       = 208'hC55072706572206F64696F207072657469756D206E65632E2046;
        inPKT[81]       = 208'hC55175736365207365642072697375732070656C6C656E746573;
        inPKT[82]       = 208'hC5527175652C20636F6E76616C6C69732073656D20656765742C;
        inPKT[83]       = 208'hC5532068656E64726572697420657261742E204D6F7262692073;
        inPKT[84]       = 208'hC5546F64616C6573207665686963756C61206C6F626F72746973;
        inPKT[85]       = 208'hC5552E2041656E65616E206120746F72746F7220637572737573;
        inPKT[86]       = 208'hC5562C207363656C65726973717565206C6967756C6120706F72;
        inPKT[87]       = 208'hC557747469746F722C20656765737461732065726F732E204475;
        inPKT[88]       = 208'hC55869732074696E636964756E7420746F72746F722069642070;
        inPKT[89]       = 208'hC5596F737565726520677261766964612E20496E20636F6E7661;
        inPKT[90]       = 208'hC55A6C6C6973206D6920696420697073756D206D616C65737561;
        inPKT[91]       = 208'hC55B64612C2075742064696374756D2065726F7320696D706572;
        inPKT[92]       = 208'hC55C646965742E2050726F696E20756C6C616D636F727065722C;
        inPKT[93]       = 208'hC55D206D61757269732069642076617269757320636F6E677565;
        inPKT[94]       = 208'hC55E2C2065726F732073617069656E2072686F6E637573206D69;
        inPKT[95]       = 208'hC55F2C20617420617563746F72206E657175652061726375206C;
        inPKT[96]       = 208'hC560616F72656574206469616D2E0D0A0D0A467573636520706F;
        inPKT[97]       = 208'hC56172747469746F72206C696265726F20617263752C206C6163;
        inPKT[98]       = 208'hC562696E69612068656E647265726974206469616D20636F6E76;
        inPKT[99]       = 208'hC563616C6C6973207365642E2050686173656C6C7573206E6F6E;
        inPKT[100]      = 208'hC564207475727069732070686172657472612C20756C6C616D63;
        inPKT[101]      = 208'hC5656F72706572206E657175652076656C2C20736F6C6C696369;
        inPKT[102]      = 208'hC566747564696E2076656C69742E2050656C6C656E7465737175;
        inPKT[103]      = 208'hC56765206861626974616E74206D6F7262692074726973746971;
        inPKT[104]      = 208'hC56875652073656E6563747573206574206E6574757320657420;
        inPKT[105]      = 208'hC5696D616C6573756164612066616D6573206163207475727069;
        inPKT[106]      = 208'hC56A7320656765737461732E204E616D206E6563207361706965;
        inPKT[107]      = 208'hC56B6E206D6F6C65737469652C2064696374756D206D61737361;
        inPKT[108]      = 208'hC56C20656765742C2065676573746173206F64696F2E20457469;
        inPKT[109]      = 208'hC56D616D20617263752073617069656E2C207072657469756D20;
        inPKT[110]      = 208'hC56E61206D6F6C6C697320612C2076756C707574617465206E6F;
        inPKT[111]      = 208'hC56F6E20657261742E205574207669746165206E696268206C6F;
        inPKT[112]      = 208'hC570626F72746973206C65637475732066617563696275732070;
        inPKT[113]      = 208'hC5716F7274612065752073697420616D6574206E69736C2E204D;
        inPKT[114]      = 208'hC5726F72626920706F72747469746F722076656C697420657520;
        inPKT[115]      = 208'hC573646F6C6F72206C616F726565742C2073697420616D657420;
        inPKT[116]      = 208'hC574696D7065726469657420656E696D20736F64616C65732E20;
        inPKT[117]      = 208'hC5754E756C6C616D20756C6C616D636F72706572207475727069;
        inPKT[118]      = 208'hC576732061742070656C6C656E74657371756520766172697573;
        inPKT[119]      = 208'hC5772E20566976616D757320657520696D70657264696574206E;
        inPKT[120]      = 208'hC578657175652E20536564207175697320617563746F7220616E;
        inPKT[121]      = 208'hC57974652E204D61757269732073656D70657220697073756D20;
        inPKT[122]      = 208'hC57A7365642064756920706F73756572652C20617420616C6971;
        inPKT[123]      = 208'hC57B75616D206D6574757320656C656966656E642E204E756C6C;
        inPKT[124]      = 208'hC57C616D2074726973746971756520656C656966656E64206572;
        inPKT[125]      = 208'hC57D6F732C2065676574206665726D656E74756D20697073756D;
        inPKT[126]      = 208'hC57E20656C656D656E74756D206E65632E0D0A0D0A50656C6C65;
        inPKT[127]      = 208'hC57F6E7465737175652068656E64726572697420626962656E64;
        inPKT[128]      = 208'hC580756D206C6967756C612C20657420736F64616C6573206D61;
        inPKT[129]      = 208'hC581676E61206461706962757320696E2E20496E20616C697175;
        inPKT[130]      = 208'hC582657420746F72746F72206567657420636F6E736563746574;
        inPKT[131]      = 208'hC583757220636F6E73656374657475722E205175697371756520;
        inPKT[132]      = 208'hC58474726973746971756520726973757320657261742C206574;
        inPKT[133]      = 208'hC58520616C697175657420656C697420616C6971756574206575;
        inPKT[134]      = 208'hC5862E20496E7465676572206E6F6E206D61676E6120696E2066;
        inPKT[135]      = 208'hC587656C697320706F72747469746F722073616769747469732E;
        inPKT[136]      = 208'hC58820517569737175652076697665727261206F726369206163;
        inPKT[137]      = 208'hC5892072757472756D206C616F726565742E2041656E65616E20;
        inPKT[138]      = 208'hC58A636F6E76616C6C69732064696374756D207475727069732C;
        inPKT[139]      = 208'hC58B2065742066696E696275732073617069656E20636F6E6775;
        inPKT[140]      = 208'hC58C6520696E2E2053656420612065726174206F726E6172652C;
        inPKT[141]      = 208'hC58D206D6F6C6C6973206E69736C2061632C206469676E697373;
        inPKT[142]      = 208'hC58E696D206E657175652E2051756973717565206D616C657375;
        inPKT[143]      = 208'hC58F61646120706F73756572652074757270697320657520756C;
        inPKT[144]      = 208'hC5906C616D636F727065722E20446F6E65632076697665727261;
        inPKT[145]      = 208'hC59120626962656E64756D206E756E632C2064696374756D2069;
        inPKT[146]      = 208'hC5926D70657264696574206E65717565206D6178696D75732069;
        inPKT[147]      = 208'hC5936E2E20446F6E656320757420756C74726963657320646F6C;
        inPKT[148]      = 208'hC5946F722E20566976616D757320736564206175677565207072;
        inPKT[149]      = 208'hC595657469756D2C20766F6C757470617420657261742061632C;
        inPKT[150]      = 208'hC59620706F727461206469616D2E204D617572697320696E2070;
        inPKT[151]      = 208'hC5977572757320756C747269636965732C207375736369706974;
        inPKT[152]      = 208'hC598206469616D207365642C2074696E636964756E7420656E69;
        inPKT[153]      = 208'hC5996D2E20446F6E6563207175697320706F7375657265206E69;
        inPKT[154]      = 208'hC59A62682E20496E206861632068616269746173736520706C61;
        inPKT[155]      = 208'hC59B7465612064696374756D73742E0D0A0D0A4D6F726269206F;
        inPKT[156]      = 208'hC59C726E617265206A7573746F206174207175616D2066617563;
        inPKT[157]      = 208'hC59D696275732C2073697420616D6574206D6F6C657374696520;
        inPKT[158]      = 208'hC59E6C656F206375727375732E204D6175726973206C616F7265;
        inPKT[159]      = 208'hC59F657420616E74652061206D65747573206566666963697475;
        inPKT[160]      = 208'hC5A072207661726975732E205365642076656C206F7263692073;
        inPKT[161]      = 208'hC5A161676974746973206E756E6320626C616E64697420636F6E;
        inPKT[162]      = 208'hC5A27365717561742E205072616573656E74206D616C65737561;
        inPKT[163]      = 208'hC5A36461206E6571756520717569732064696374756D20646967;
        inPKT[164]      = 208'hC5A46E697373696D2E20446F6E656320666163696C6973697320;
        inPKT[165]      = 208'hC5A573697420616D65742076656C6974206575206C6F626F7274;
        inPKT[166]      = 208'hC5A669732E204E756C6C616D20626C616E64697420656C656D65;
        inPKT[167]      = 208'hC5A76E74756D206D61757269732C20766974616520656C656D65;
        inPKT[168]      = 208'hC5A86E74756D20646F6C6F722068656E64726572697420766974;
        inPKT[169]      = 208'hC5A961652E204675736365206D6F6C65737469652C20656C6974;
        inPKT[170]      = 208'hC5AA20757420616C697175657420766F6C75747061742C206E65;
        inPKT[171]      = 208'hC5AB7175652076656C6974207072657469756D2061756775652C;
        inPKT[172]      = 208'hC5AC206672696E67696C6C6120636F6E64696D656E74756D206A;
        inPKT[173]      = 208'hC5AD7573746F2073617069656E2061206A7573746F2E20506861;
        inPKT[174]      = 208'hC5AE73656C6C7573207175697320617563746F72206C6F72656D;
        inPKT[175]      = 208'hC5AF2C20696E20616C697175616D206E756E632E20557420656C;
        inPKT[176]      = 208'hC5B0656966656E6420616E7465206574206E697369206D6F6C65;
        inPKT[177]      = 208'hC5B17374696520636F6E76616C6C69732069642065742073656D;
        inPKT[178]      = 208'hC5B22E2053656420616320626962656E64756D20617263752E20;
        inPKT[179]      = 208'hC5B3467573636520766573746962756C756D206E756E63206567;
        inPKT[180]      = 208'hC5B465742074656C6C7573206665726D656E74756D2C206E6563;
        inPKT[181]      = 208'hC5B52072686F6E637573206D6173736120636F6D6D6F646F2E20;
        inPKT[182]      = 208'hC5B64D616563656E6173206964206E756E63206E6F6E20657820;
        inPKT[183]      = 208'hC5B7766573746962756C756D206F726E617265207574206E6563;
        inPKT[184]      = 208'hC5B82065726F732E20416C697175616D20656666696369747572;
        inPKT[185]      = 208'hC5B920636F6D6D6F646F206469616D206964206C6F626F727469;
        inPKT[186]      = 208'hC5BA732E205365642061632074656D706F72206C65637475732E;
        inPKT[187]      = 208'hC5BB204E756E6320656C656D656E74756D207574206C65637475;
        inPKT[188]      = 208'hC5BC732061632074696E636964756E742E20557420696163756C;
        inPKT[189]      = 208'hC5BD6973206E756C6C61207175697320657820656C656D656E74;
        inPKT[190]      = 208'hC5BE756D2C20616C69717565742073656D706572206D61676E61;
        inPKT[191]      = 208'hC5BF20656C656966656E642E0D0A0D0A43757261626974757220;
        inPKT[192]      = 208'hC5C0746F72746F72206E69736C2C20756C747269636965732069;
        inPKT[193]      = 208'hC5C16E206E657175652061632C20616363756D73616E20636F6E;
        inPKT[194]      = 208'hC5C2736571756174206D657475732E204D616563656E6173206D;
        inPKT[195]      = 208'hC5C3617373612073617069656E2C206D617474697320696E2076;
        inPKT[196]      = 208'hC5C4656E656E617469732073697420616D65742C20617563746F;
        inPKT[197]      = 208'hC5C5722073697420616D657420656E696D2E204E756E63207669;
        inPKT[198]      = 208'hC5C6746165206D6574757320636F6D6D6F646F2C206D61747469;
        inPKT[199]      = 208'hC5C773206D617373612073697420616D65742C20766172697573;
        inPKT[200]      = 208'hC5C8206C6F72656D2E204E756E6320696E20656C697420656C69;
        inPKT[201]      = 208'hC5C9742E204E756E63206F726E61726520636F6E736563746574;
        inPKT[202]      = 208'hC5CA7572206D61676E612C2073697420616D657420706F727474;
        inPKT[203]      = 208'hC5CB69746F7220617263752072686F6E6375732065752E205375;
        inPKT[204]      = 208'hC5CC7370656E6469737365207363656C6572697371756520756C;
        inPKT[205]      = 208'hC5CD74726963696573206578206120616C697175616D2E205375;
        inPKT[206]      = 208'hC5CE7370656E64697373652072757472756D20736F6C6C696369;
        inPKT[207]      = 208'hC5CF747564696E206E756E632C206E6F6E20636F6E76616C6C69;
        inPKT[208]      = 208'hC5D07320747572706973206C616F726565742073697420616D65;
        inPKT[209]      = 208'hC5D1742E2041656E65616E20612066696E69627573206D617572;
        inPKT[210]      = 208'hC5D269732C207175697320637572737573206E756E632E20496E;
        inPKT[211]      = 208'hC5D32066657567696174206475692076656C2075726E61207365;
        inPKT[212]      = 208'hC5D46D7065722066617563696275732E204D617572697320756C;
        inPKT[213]      = 208'hC5D5747269636965732061742074757270697320656765742070;
        inPKT[214]      = 208'hC5D6656C6C656E7465737175652E205072616573656E74207369;
        inPKT[215]      = 208'hC5D77420616D6574206C6967756C6120636F6E76616C6C69732C;
        inPKT[216]      = 208'hC5D820656C656D656E74756D206E756C6C6120756C6C616D636F;
        inPKT[217]      = 208'hC5D9727065722C20616C697175616D2075726E612E2045746961;
        inPKT[218]      = 208'hC5DA6D207175616D20656C69742C20706F737565726520757420;
        inPKT[219]      = 208'hC5DB7175616D20656765742C2066696E6962757320736F6C6C69;
        inPKT[220]      = 208'hC5DC6369747564696E206E756C6C612E20496E20737573636970;
        inPKT[221]      = 208'hC5DD697420656E696D2065742065726F732066696E696275732C;
        inPKT[222]      = 208'hC5DE207574207363656C657269737175652074656C6C75732066;
        inPKT[223]      = 208'hC5DF6575676961742E20437572616269747572206E6F6E206D61;
        inPKT[224]      = 208'hC5E07373612076617269757320646F6C6F722067726176696461;
        inPKT[225]      = 208'hC5E120656C656D656E74756D20717569732075742066656C6973;
        inPKT[226]      = 208'hC5E22E2050686173656C6C757320657569736D6F642069707375;
        inPKT[227]      = 208'hC5E36D20656765742076656C6974206C6F626F727469732C2065;
        inPKT[228]      = 208'hC5E467657420706F727461206D61757269732074656D7075732E;
        inPKT[229]      = 208'hC5E52053656420696D7065726469657420766F6C757470617420;
        inPKT[230]      = 208'hC5E674656C6C75732065752074696E636964756E742E0D0A0D0A;
        inPKT[231]      = 208'hC5E755742076656C206D69206174206D65747573206672696E67;
        inPKT[232]      = 208'hC5E8696C6C6120677261766964612E205072616573656E742065;
        inPKT[233]      = 208'hC5E9726F73206E6962682C206375727375732065676573746173;
        inPKT[234]      = 208'hC5EA2074696E636964756E7420736F64616C65732C207363656C;
        inPKT[235]      = 208'hC5EB65726973717565206E65632066656C69732E20496E746567;
        inPKT[236]      = 208'hC5EC657220696D70657264696574206D616C657375616461206E;
        inPKT[237]      = 208'hC5ED69736C20616C69717565742076656E656E617469732E2049;
        inPKT[238]      = 208'hC5EE6E74656765722073656420706F72747469746F7220697073;
        inPKT[239]      = 208'hC5EF756D2E20496E746567657220636F6D6D6F646F2066657567;
        inPKT[240]      = 208'hC5F069617420746F72746F722C206575206C6F626F7274697320;
        inPKT[241]      = 208'hC5F1617567756520656C656D656E74756D2073697420616D6574;
        inPKT[242]      = 208'hC5F22E20446F6E656320766573746962756C756D206C6967756C;
        inPKT[243]      = 208'hC5F3612061756775652C2065742066696E696275732061726375;
        inPKT[244]      = 208'hC5F420706F72746120696E2E204E756C6C612073656D2074656C;
        inPKT[245]      = 208'hC5F56C75732C20756C6C616D636F727065722061742063757273;
        inPKT[246]      = 208'hC5F6757320612C20706F7274612073697420616D6574206D6167;
        inPKT[247]      = 208'hC5F76E612E204E756E6320766974616520696D70657264696574;
        inPKT[248]      = 208'hC5F82070757275732C206E656320736F6C6C696369747564696E;
        inPKT[249]      = 208'hC5F92074656C6C75732E20416C697175616D206572617420766F;
        inPKT[250]      = 208'hC5FA6C75747061742E20536564206964206D61676E6120636F6D;
        inPKT[251]      = 208'hC5FB6D6F646F2C206C75637475732076656C697420717569732C;
        inPKT[252]      = 208'hC5FC20657569736D6F6420656E696D2E20496E7465676572206D;
        inPKT[253]      = 208'hC5FD617474697320736F64616C6573206665726D656E74756D2E;
        inPKT[254]      = 208'hC5FE205175697371756520736564206672696E67696C6C61206C;
        inPKT[255]      = 208'hC5FF6F72656D2E2043726173207665686963756C612074656D70;
        inPKT[256]      = 208'hC50075732073617069656E20757420636F6E6775652E20447569;
        inPKT[257]      = 208'hC501732073617069656E20656E696D2C20706F727461206E6563;
        inPKT[258]      = 208'hC502206C656F2069642C2065666669636974757220706F737565;
        inPKT[259]      = 208'hC5037265206C696265726F2E204E756C6C616D2061632074656D;
        inPKT[260]      = 208'hC504706F72206D657475732E205365642076656C207475727069;
        inPKT[261]      = 208'hC5057320666575676961742C20696163756C6973206175677565;
        inPKT[262]      = 208'hC50620717569732C2074696E636964756E74207475727069732E;
        inPKT[263]      = 208'hC5070D0A0D0A566976616D757320706F737565726520706F7274;
        inPKT[264]      = 208'hC5087469746F722061756775652C207661726975732061636375;
        inPKT[265]      = 208'hC5096D73616E20656C69742076756C7075746174652065676574;
        inPKT[266]      = 208'hC50A2E205175697371756520736564206D616C65737561646120;
        inPKT[267]      = 208'hC50B6E69736C2E20496E74657264756D206574206D616C657375;
        inPKT[268]      = 208'hC50C6164612066616D657320616320616E746520697073756D20;
        inPKT[269]      = 208'hC50D7072696D697320696E2066617563696275732E204E756E63;
        inPKT[270]      = 208'hC50E20747572706973206469616D2C2073757363697069742061;
        inPKT[271]      = 208'hC50F632065726F732076656C2C2074656D7075732076656E656E;
        inPKT[272]      = 208'hC5106174697320697073756D2E2044756973206C756374757320;
        inPKT[273]      = 208'hC51172686F6E637573206D617373612E20467573636520757420;
        inPKT[274]      = 208'hC5126C6163696E6961207475727069732E20566976616D757320;
        inPKT[275]      = 208'hC51372757472756D2074656C6C75732061756775652C20617420;
        inPKT[276]      = 208'hC5146F726E617265206E69736C20666163696C69736973206574;
        inPKT[277]      = 208'hC5152E204E756E6320736564206E6973692072697375732E2049;
        inPKT[278]      = 208'hC5166E746567657220656C656D656E74756D206D617572697320;
        inPKT[279]      = 208'hC5177175616D2C207574207665686963756C61206D6175726973;
        inPKT[280]      = 208'hC51820636F6E6775652065752E0D0A0D0A467573636520612074;
        inPKT[281]      = 208'hC519656C6C75732073697420616D65742065726174206665726D;
        inPKT[282]      = 208'hC51A656E74756D207363656C657269737175652E204375726162;
        inPKT[283]      = 208'hC51B6974757220696E2076656C697420617420656E696D206C61;
        inPKT[284]      = 208'hC51C63696E6961207665686963756C61206163206964206A7573;
        inPKT[285]      = 208'hC51D746F2E2050726F696E206E6F6E20646F6C6F722065666669;
        inPKT[286]      = 208'hC51E63697475722C2074696E636964756E74206F64696F206575;
        inPKT[287]      = 208'hC51F2C20666175636962757320656E696D2E2050656C6C656E74;
        inPKT[288]      = 208'hC52065737175652064617069627573206F726369206163206C6F;
        inPKT[289]      = 208'hC52172656D20696163756C69732C2073697420616D657420626C;
        inPKT[290]      = 208'hC522616E6469742061726375207472697374697175652E204165;
        inPKT[291]      = 208'hC5236E65616E2074726973746971756520746F72746F72206E65;
        inPKT[292]      = 208'hC52463206A7573746F20616C697175616D2C20696E2070726574;
        inPKT[293]      = 208'hC52569756D2066656C6973206D6F6C65737469652E2053656420;
        inPKT[294]      = 208'hC52665742074656D7075732061756775652E204E756C6C612066;
        inPKT[295]      = 208'hC52772696E67696C6C6120656C656966656E6420697073756D20;
        inPKT[296]      = 208'hC52876697665727261206375727375732E20416C697175616D20;
        inPKT[297]      = 208'hC5296D6178696D7573206665726D656E74756D206E6962682061;
        inPKT[298]      = 208'hC52A6320616363756D73616E2E204E756C6C6120666163696C69;
        inPKT[299]      = 208'hC52B73692E20566573746962756C756D20666163696C69736973;
        inPKT[300]      = 208'hC52C206C656F20656765737461732073656D206D617474697320;
        inPKT[301]      = 208'hC52D636F6E6775652E204D617572697320766974616520657820;
        inPKT[302]      = 208'hC52E6174207269737573206461706962757320656C656966656E;
        inPKT[303]      = 208'hC52F642E20496E74656765722075742065726F7320636F6E6775;
        inPKT[304]      = 208'hC530652C20706F72747469746F7220616E7465206E6F6E2C2069;
        inPKT[305]      = 208'hC5316E74657264756D20646F6C6F722E0D0A0D0A566573746962;
        inPKT[306]      = 208'hC532756C756D20656C656966656E64206D617572697320657520;
        inPKT[307]      = 208'hC5336E6973692064696374756D20677261766964612E20447569;
        inPKT[308]      = 208'hC53473206D6F6C6C6973206469616D2076656C20656E696D2074;
        inPKT[309]      = 208'hC535656D7075732C2076697461652064617069627573206D6173;
        inPKT[310]      = 208'hC53673612073616769747469732E204E756C6C61207574206175;
        inPKT[311]      = 208'hC53763746F7220746F72746F722E204D6F72626920736564206C;
        inPKT[312]      = 208'hC5386F72656D2075726E612E204675736365206D61747469732C;
        inPKT[313]      = 208'hC539206D61676E6120616320636F6E64696D656E74756D206665;
        inPKT[314]      = 208'hC53A75676961742C206D6173736120647569206D6178696D7573;
        inPKT[315]      = 208'hC53B206E756C6C612C20657520616C6971756574206E65717565;
        inPKT[316]      = 208'hC53C206D6175726973206120657261742E205175697371756520;
        inPKT[317]      = 208'hC53D617563746F722065737420757420696E74657264756D2063;
        inPKT[318]      = 208'hC53E6F6E73656374657475722E20446F6E656320656765742064;
        inPKT[319]      = 208'hC53F69676E697373696D20746F72746F722C2068656E64726572;
        inPKT[320]      = 208'hC5406974206D617474697320657261742E2050656C6C656E7465;
        inPKT[321]      = 208'hC54173717565206861626974616E74206D6F7262692074726973;
        inPKT[322]      = 208'hC54274697175652073656E6563747573206574206E6574757320;
        inPKT[323]      = 208'hC5436574206D616C6573756164612066616D6573206163207475;
        inPKT[324]      = 208'hC5447270697320656765737461732E2051756973717565206F72;
        inPKT[325]      = 208'hC5456E617265207661726975732074656D7075732E0D0A0D0A4D;
        inPKT[326]      = 208'hC5466F7262692072757472756D20616E7465206E6962682C2061;
        inPKT[327]      = 208'hC5472076697665727261206E756C6C612068656E647265726974;
        inPKT[328]      = 208'hC54820696E2E2050726F696E2073757363697069742065676573;
        inPKT[329]      = 208'hC54974617320657261742C20757420617563746F72206F726369;
        inPKT[330]      = 208'hC54A206D617474697320612E2050656C6C656E74657371756520;
        inPKT[331]      = 208'hC54B6C7563747573206672696E67696C6C6120656C6974207574;
        inPKT[332]      = 208'hC54C206C6163696E69612E205574206574206D61737361206E75;
        inPKT[333]      = 208'hC54D6C6C612E20536564206174206672696E67696C6C61206C6F;
        inPKT[334]      = 208'hC54E72656D2E2050726F696E206772617669646120616363756D;
        inPKT[335]      = 208'hC54F73616E2072697375732073656420626962656E64756D2E20;
        inPKT[336]      = 208'hC5504D616563656E6173206D616C657375616461206F64696F20;
        inPKT[337]      = 208'hC55175742076656C697420657569736D6F642064617069627573;
        inPKT[338]      = 208'hC5522E0D0A0D0A457469616D20636F6E677565206D6174746973;
        inPKT[339]      = 208'hC55320696163756C69732E204D61757269732076697461652065;
        inPKT[340]      = 208'hC55466666963697475722073656D2E205365642070756C76696E;
        inPKT[341]      = 208'hC555617220646F6C6F72207574206D6920657569736D6F642068;
        inPKT[342]      = 208'hC556656E6472657269742E204E756C6C616D2061742067726176;
        inPKT[343]      = 208'hC55769646120646F6C6F722E204D6F726269206C656F20747572;
        inPKT[344]      = 208'hC5587069732C20636F6E677565206E656320616C697175616D20;
        inPKT[345]      = 208'hC55975742C20636F6D6D6F646F20696E206E756E632E204E756C;
        inPKT[346]      = 208'hC55A6C61206174206661756369627573206C656F2C2065752066;
        inPKT[347]      = 208'hC55B657567696174206C616375732E204675736365206E6F6E20;
        inPKT[348]      = 208'hC55C65676573746173207475727069732E205175697371756520;
        inPKT[349]      = 208'hC55D766974616520697073756D206D692E204E756E63206E6F6E;
        inPKT[350]      = 208'hC55E206F7263692073697420616D6574206E6973692076617269;
        inPKT[351]      = 208'hC55F757320706F72747469746F7220696E2076756C7075746174;
        inPKT[352]      = 208'hC5606520746F72746F722E204E756E6320636F6E76616C6C6973;
        inPKT[353]      = 208'hC5612067726176696461206469616D206120756C747269636965;
        inPKT[354]      = 208'hC562732E2051756973717565206575206A7573746F20636F6E64;
        inPKT[355]      = 208'hC563696D656E74756D2C20766172697573206469616D2076656C;
        inPKT[356]      = 208'hC5642C20766573746962756C756D206D617373612E0D0A0D0A50;
        inPKT[357]      = 208'hC565656C6C656E7465737175652070656C6C656E746573717565;
        inPKT[358]      = 208'hC5662073617069656E206E657175652C20617563746F72206D61;
        inPKT[359]      = 208'hC5676C65737561646120657261742068656E647265726974206E;
        inPKT[360]      = 208'hC56865632E204E756C6C6120706C616365726174206469616D20;
        inPKT[361]      = 208'hC56968656E647265726974206D6173736120626962656E64756D;
        inPKT[362]      = 208'hC56A2C2061206D6F6C65737469652066656C69732068656E6472;
        inPKT[363]      = 208'hC56B657269742E204D617572697320657569736D6F642076656E;
        inPKT[364]      = 208'hC56C656E61746973206A7573746F2C20757420617563746F7220;
        inPKT[365]      = 208'hC56D656C697420616C69717565742075742E2046757363652061;
        inPKT[366]      = 208'hC56E6C69717565742C207175616D207574206469676E69737369;
        inPKT[367]      = 208'hC56F6D2068656E6472657269742C206D61757269732074757270;
        inPKT[368]      = 208'hC5706973206469676E697373696D20746F72746F722C20656765;
        inPKT[369]      = 208'hC571742070656C6C656E7465737175652076656C6974206F7263;
        inPKT[370]      = 208'hC57269206E6563207175616D2E204E756E632065676573746173;
        inPKT[371]      = 208'hC5732070656C6C656E7465737175652072697375732E20437572;
        inPKT[372]      = 208'hC5746162697475722073757363697069742074656D707573206C;
        inPKT[373]      = 208'hC575616375732C2065676574207072657469756D20656C697420;
        inPKT[374]      = 208'hC57674696E636964756E74206E6F6E2E20437261732075726E61;
        inPKT[375]      = 208'hC577206C6F72656D2C20706C61636572617420766F6C75747061;
        inPKT[376]      = 208'hC5787420696D706572646965742073697420616D65742C206567;
        inPKT[377]      = 208'hC57965737461732076656C206F7263692E0D0A0D0A50656C6C65;
        inPKT[378]      = 208'hC57A6E74657371756520736F64616C6573206665726D656E7475;
        inPKT[379]      = 208'hC57B6D206E69736C2C206174206672696E67696C6C6120647569;
        inPKT[380]      = 208'hC57C2073656D706572206665726D656E74756D2E204E756C6C61;
        inPKT[381]      = 208'hC57D6D20706C6163657261742076656C206D692068656E647265;
        inPKT[382]      = 208'hC57E72697420656C656D656E74756D2E20457469616D206E6F6E;
        inPKT[383]      = 208'hC57F20697073756D2065782E204E616D206163207363656C6572;
        inPKT[384]      = 208'hC5806973717565206E6962682C2076656C20666163696C697369;
        inPKT[385]      = 208'hC58173206D692E20446F6E65632065676573746173206C616F72;
        inPKT[386]      = 208'hC5826565742065726F732C206567657420766F6C757470617420;
        inPKT[387]      = 208'hC5836D657475732E205072616573656E7420616363756D73616E;
        inPKT[388]      = 208'hC58420626962656E64756D206E69736C206E65632076656E656E;
        inPKT[389]      = 208'hC585617469732E205365642072757472756D206D692061207375;
        inPKT[390]      = 208'hC5867363697069742070686172657472612E2053656420736974;
        inPKT[391]      = 208'hC58720616D657420696E74657264756D207475727069732E2041;
        inPKT[392]      = 208'hC5886C697175616D206575206E69626820746F72746F722E2044;
        inPKT[393]      = 208'hC5896F6E65632066617563696275732064617069627573206E69;
        inPKT[394]      = 208'hC58A73692C20736564206C616F72656574206F72636920736365;
        inPKT[395]      = 208'hC58B6C6572697371756520696E2E0D0A0D0A4D61757269732069;
        inPKT[396]      = 208'hC58C6E2066656C6973206665726D656E74756D2C20636F6E7661;
        inPKT[397]      = 208'hC58D6C6C69732061756775652076656C2C20706F737565726520;
        inPKT[398]      = 208'hC58E6D692E2050656C6C656E746573717565207363656C657269;
        inPKT[399]      = 208'hC58F737175652072686F6E637573206A7573746F2C2065752070;
        inPKT[400]      = 208'hC590756C76696E617220656E696D2070756C76696E6172207665;
        inPKT[401]      = 208'hC5916C2E204D616563656E6173207068617265747261206C6962;
        inPKT[402]      = 208'hC59265726F206D61676E612C20616320736F6C6C696369747564;
        inPKT[403]      = 208'hC593696E206C656F206D6F6C6C6973206E6F6E2E204E756C6C61;
        inPKT[404]      = 208'hC59420656C656D656E74756D206F726E61726520656765737461;
        inPKT[405]      = 208'hC595732E20436C61737320617074656E74207461636974692073;
        inPKT[406]      = 208'hC5966F63696F737175206164206C69746F726120746F72717565;
        inPKT[407]      = 208'hC5976E742070657220636F6E75626961206E6F737472612C2070;
        inPKT[408]      = 208'hC598657220696E636570746F732068696D656E61656F732E2050;
        inPKT[409]      = 208'hC59972616573656E74206175677565206D61757269732C207268;
        inPKT[410]      = 208'hC59A6F6E637573207175697320657374206E6F6E2C206D6F6C6C;
        inPKT[411]      = 208'hC59B697320636F6E76616C6C69732066656C69732E2053757370;
        inPKT[412]      = 208'hC59C656E646973736520666163696C697369732C206F72636920;
        inPKT[413]      = 208'hC59D7669746165206C6163696E69612074656D706F722C206C65;
        inPKT[414]      = 208'hC59E637475732073617069656E206D6174746973207269737573;
        inPKT[415]      = 208'hC59F2C206E6F6E20736167697474697320656C6974206E657175;
        inPKT[416]      = 208'hC5A0652071756973206A7573746F2E20446F6E6563206D616C65;
        inPKT[417]      = 208'hC5A17375616461206C6163696E6961206475692E205068617365;
        inPKT[418]      = 208'hC5A26C6C75732068656E647265726974206D6175726973206D61;
        inPKT[419]      = 208'hC5A3757269732C20736564206672696E67696C6C61206C696265;
        inPKT[420]      = 208'hC5A4726F206672696E67696C6C6120696E2E2053656420617420;
        inPKT[421]      = 208'hC5A56C6967756C6120696E206A7573746F2066696E6962757320;
        inPKT[422]      = 208'hC5A676756C7075746174652E204E756E6320637572737573206E;
        inPKT[423]      = 208'hC5A7657175652073697420616D657420617263752074696E6369;
        inPKT[424]      = 208'hC5A864756E742C2076697461652070686172657472612073656D;
        inPKT[425]      = 208'hC5A920706F72747469746F722E20416C697175616D206D617474;
        inPKT[426]      = 208'hC5AA69732C206A7573746F206E6F6E20657569736D6F6420636F;
        inPKT[427]      = 208'hC5AB6E76616C6C69732C206E756E63206D6920636F6E73657175;
        inPKT[428]      = 208'hC5AC6174206573742C206E656320736F6C6C696369747564696E;
        inPKT[429]      = 208'hC5AD206C65637475732073617069656E2076656C206F64696F2E;
        inPKT[430]      = 208'hC5AE20496E2074656D706F72206572617420646F6C6F722C2073;
        inPKT[431]      = 208'hC5AF6564207665686963756C612075726E6120636F6E73657175;
        inPKT[432]      = 208'hC5B06174207365642E0D0A0D0A4E616D2072686F6E6375732069;
        inPKT[433]      = 208'hC5B164206D6175726973206E6563206469676E697373696D2E20;
        inPKT[434]      = 208'hC5B2496E20696D7065726469657420756C747269636573206572;
        inPKT[435]      = 208'hC5B36174206E656320736F6C6C696369747564696E2E20496E74;
        inPKT[436]      = 208'hC5B4656765722073656420636F6E64696D656E74756D2065726F;
        inPKT[437]      = 208'hC5B5732E20446F6E65632065676574206E756E63206964206D61;
        inPKT[438]      = 208'hC5B6757269732074726973746971756520706F72747469746F72;
        inPKT[439]      = 208'hC5B7206C616F72656574207669746165206D657475732E204E75;
        inPKT[440]      = 208'hC5B86C6C6120666163696C6973692E204E756C6C616D20657520;
        inPKT[441]      = 208'hC5B96C616375732061206469616D207472697374697175652065;
        inPKT[442]      = 208'hC5BA676573746173206E6F6E20696163756C6973206D65747573;
        inPKT[443]      = 208'hC5BB2E20416C697175616D20696E2074656D706F722065726174;
        inPKT[444]      = 208'hC5BC2C20696420636F6E677565206D617373612E20566976616D;
        inPKT[445]      = 208'hC5BD75732076656C20746F72746F72207669746165206E696268;
        inPKT[446]      = 208'hC5BE20636F6D6D6F646F206C6F626F7274697320717569732061;
        inPKT[447]      = 208'hC5BF20697073756D2E2050726F696E20766F6C75747061742071;
        inPKT[448]      = 208'hC5C075616D206E6F6E2066656C69732074656D7075732C206964;
        inPKT[449]      = 208'hC5C120706F737565726520646F6C6F722074656D706F722E2050;
        inPKT[450]      = 208'hC5C272616573656E742076697461652074696E636964756E7420;
        inPKT[451]      = 208'hC5C373617069656E2E204D616563656E617320666163696C6973;
        inPKT[452]      = 208'hC5C46973206D617474697320616E746520717569732076617269;
        inPKT[453]      = 208'hC5C575732E20446F6E65632070656C6C656E7465737175652065;
        inPKT[454]      = 208'hC5C6726F7320666575676961742074696E636964756E7420636F;
        inPKT[455]      = 208'hC5C76E64696D656E74756D2E2050726F696E2066617563696275;
        inPKT[456]      = 208'hC5C87320766F6C7574706174206D692073656420736167697474;
        inPKT[457]      = 208'hC5C969732E0D0A0D0A44756973206772617669646120656C656D;
        inPKT[458]      = 208'hC5CA656E74756D20696E74657264756D2E2050726F696E207369;
        inPKT[459]      = 208'hC5CB7420616D6574207175616D206C6967756C612E2050686173;
        inPKT[460]      = 208'hC5CC656C6C757320636F6D6D6F646F2C2075726E6120696E2063;
        inPKT[461]      = 208'hC5CD6F6E67756520766F6C75747061742C206C6967756C612065;
        inPKT[462]      = 208'hC5CE78207068617265747261206C6967756C612C20696E206469;
        inPKT[463]      = 208'hC5CF6374756D206D61676E61206F726369206E6563206D617572;
        inPKT[464]      = 208'hC5D069732E204E756E6320617563746F7220636F6E7365637465;
        inPKT[465]      = 208'hC5D174757220766F6C75747061742E204D6F7262692074696E63;
        inPKT[466]      = 208'hC5D26964756E74206E69626820757420656E696D206566666963;
        inPKT[467]      = 208'hC5D36974757220677261766964612E2043757261626974757220;
        inPKT[468]      = 208'hC5D47669746165207175616D2065726F732E2044756973206672;
        inPKT[469]      = 208'hC5D5696E67696C6C6120616320746F72746F7220696E2074696E;
        inPKT[470]      = 208'hC5D6636964756E742E204E756E632076656C206D617572697320;
        inPKT[471]      = 208'hC5D772697375732E20446F6E656320656C656966656E64206C69;
        inPKT[472]      = 208'hC5D867756C61207361676974746973206E6973692066696E6962;
        inPKT[473]      = 208'hC5D975732C2061207363656C65726973717565206C696265726F;
        inPKT[474]      = 208'hC5DA2070656C6C656E7465737175652E20566573746962756C75;
        inPKT[475]      = 208'hC5DB6D20747269737469717565206D61737361206E6962682C20;
        inPKT[476]      = 208'hC5DC617420766573746962756C756D206D61676E612066696E69;
        inPKT[477]      = 208'hC5DD6275732065752E0D0A0D0A43757261626974757220696D70;
        inPKT[478]      = 208'hC5DE6572646965742070757275732065676574206E756E632075;
        inPKT[479]      = 208'hC5DF6C7472696365732C2076697461652076656E656E61746973;
        inPKT[480]      = 208'hC5E0206D6173736120636F6D6D6F646F2E2050656C6C656E7465;
        inPKT[481]      = 208'hC5E173717565206861626974616E74206D6F7262692074726973;
        inPKT[482]      = 208'hC5E274697175652073656E6563747573206574206E6574757320;
        inPKT[483]      = 208'hC5E36574206D616C6573756164612066616D6573206163207475;
        inPKT[484]      = 208'hC5E47270697320656765737461732E20496E206665726D656E74;
        inPKT[485]      = 208'hC5E5756D2061742075726E61206E6F6E20636F6E76616C6C6973;
        inPKT[486]      = 208'hC5E62E20446F6E6563206163206175677565206A7573746F2E20;
        inPKT[487]      = 208'hC5E7496E20617420656C69742065742061726375206D6178696D;
        inPKT[488]      = 208'hC5E87573206C75637475732E20467573636520657569736D6F64;
        inPKT[489]      = 208'hC5E9206E756E63206E65632076656E656E617469732061756374;
        inPKT[490]      = 208'hC5EA6F722E204C6F72656D20697073756D20646F6C6F72207369;
        inPKT[491]      = 208'hC5EB7420616D65742C20636F6E73656374657475722061646970;
        inPKT[492]      = 208'hC5EC697363696E6720656C69742E20446F6E6563206469637475;
        inPKT[493]      = 208'hC5ED6D2074656D706F722072757472756D2E2053656420656C65;
        inPKT[494]      = 208'hC5EE6966656E64206469616D206964206D6173736120696D7065;
        inPKT[495]      = 208'hC5EF72646965742C206163206F726E617265206C696265726F20;
        inPKT[496]      = 208'hC5F0656C656966656E642E204D616563656E6173206F726E6172;
        inPKT[497]      = 208'hC5F165206D65747573206E756C6C612C2073697420616D657420;
        inPKT[498]      = 208'hC5F26665726D656E74756D20656C697420616C697175616D2069;
        inPKT[499]      = 208'hC5F3642E20446F6E656320756C74726963657320746F72746F72;
        inPKT[500]      = 208'hC5F420617420616E74652068656E6472657269742C2065752073;
        inPKT[501]      = 208'hC5F561676974746973206A7573746F20756C7472696365732E0D;
        inPKT[502]      = 208'hC5F60A0D0A5072616573656E74206C7563747573207072657469;
        inPKT[503]      = 208'hC5F7756D206E657175652C2073697420616D65742070656C6C65;
        inPKT[504]      = 208'hC5F86E746573717565206D617572697320656C656D656E74756D;
        inPKT[505]      = 208'hC5F9206E6F6E2E20557420626C616E6469742070686172657472;
        inPKT[506]      = 208'hC5FA61206F64696F206E6F6E20657569736D6F642E2051756973;
        inPKT[507]      = 208'hC5FB717565207669746165206C656F20616C697175616D2C2073;
        inPKT[508]      = 208'hC5FC6F64616C65732074656C6C75732069642C20696163756C69;
        inPKT[509]      = 208'hC5FD73206D61757269732E204E616D2065666669636974757220;
        inPKT[510]      = 208'hC5FE696E2070757275732073656420616363756D73616E2E204D;
        inPKT[511]      = 208'hC5FF616563656E61732073697420616D65742063757273757320;
        inPKT[512]      = 208'hC50066656C69732E20517569737175652066617563696275732C;
        inPKT[513]      = 208'hC5012064756920657420617563746F72206C75637475732C2061;
        inPKT[514]      = 208'hC5026E7465206572617420706F73756572652065726F732C2075;
        inPKT[515]      = 208'hC5037420636F6E76616C6C6973206D65747573206C6563747573;
        inPKT[516]      = 208'hC504207669746165206C656F2E2053757370656E646973736520;
        inPKT[517]      = 208'hC505706F74656E74692E204372617320657420646F6C6F72206E;
        inPKT[518]      = 208'hC5066F6E2075726E61207363656C657269737175652074726973;
        inPKT[519]      = 208'hC50774697175652E20437261732072757472756D206E65632076;
        inPKT[520]      = 208'hC508656C69742061632073616769747469732E20446F6E656320;
        inPKT[521]      = 208'hC509656C656966656E642C206C61637573207365642067726176;
        inPKT[522]      = 208'hC50A696461206D616C6573756164612C20657820616E74652070;
        inPKT[523]      = 208'hC50B6C616365726174206C65637475732C206567657420636F6E;
        inPKT[524]      = 208'hC50C677565206D61737361206D65747573206964206C61637573;
        inPKT[525]      = 208'hC50D2E2053757370656E64697373652069642072757472756D20;
        inPKT[526]      = 208'hC50E6C65637475732E204675736365206D6178696D7573207365;
        inPKT[527]      = 208'hC50F64206C6967756C612073656420766976657272612E204E61;
        inPKT[528]      = 208'hC5106D206C7563747573206469616D20616E74652C2076697461;
        inPKT[529]      = 208'hC51165206F726E617265206E6571756520766172697573206567;
        inPKT[530]      = 208'hC51265742E0D0A0D0A50656C6C656E7465737175652061742065;
        inPKT[531]      = 208'hC5136C6974206E6962682E20566573746962756C756D20616E74;
        inPKT[532]      = 208'hC5146520697073756D207072696D697320696E20666175636962;
        inPKT[533]      = 208'hC5157573206F726369206C756374757320657420756C74726963;
        inPKT[534]      = 208'hC516657320706F737565726520637562696C6961204375726165;
        inPKT[535]      = 208'hC5173B2043757261626974757220666175636962757320646961;
        inPKT[536]      = 208'hC5186D206C656F2C206E656320657569736D6F642073656D2065;
        inPKT[537]      = 208'hC51966666963697475722075742E205574207665686963756C61;
        inPKT[538]      = 208'hC51A206175677565206163206C696265726F20696163756C6973;
        inPKT[539]      = 208'hC51B2C206E656320656C656966656E6420657820706F7274612E;
        inPKT[540]      = 208'hC51C204D6F7262692068656E6472657269742067726176696461;
        inPKT[541]      = 208'hC51D2074696E636964756E742E205072616573656E7420646F6C;
        inPKT[542]      = 208'hC51E6F72206C616375732C2074656D707573206575206672696E;
        inPKT[543]      = 208'hC51F67696C6C612073697420616D65742C20656C656966656E64;
        inPKT[544]      = 208'hC52020696E206E756C6C612E204E756C6C61206D6F6C6C697320;
        inPKT[545]      = 208'hC52165676574206D61676E61206E65632068656E647265726974;
        inPKT[546]      = 208'hC5222E20416C697175616D20636F6E76616C6C69732073656D20;
        inPKT[547]      = 208'hC52376697461652073617069656E2064696374756D2C20757420;
        inPKT[548]      = 208'hC524766573746962756C756D206C6F72656D206672696E67696C;
        inPKT[549]      = 208'hC5256C612E20446F6E65632074656C6C7573206C696265726F2C;
        inPKT[550]      = 208'hC52620666575676961742075742066696E69627573206E65632C;
        inPKT[551]      = 208'hC52720616C697175616D2073697420616D6574206F7263692E20;
        inPKT[552]      = 208'hC5284E756E63207375736369706974206E69736C206574206F72;
        inPKT[553]      = 208'hC5296E61726520766573746962756C756D2E204E756C6C616D20;
        inPKT[554]      = 208'hC52A6C6F626F727469732073617069656E206A7573746F2C2073;
        inPKT[555]      = 208'hC52B697420616D6574206469676E697373696D206E756C6C6120;
        inPKT[556]      = 208'hC52C636F6E64696D656E74756D20696E2E20536564206D6F6C65;
        inPKT[557]      = 208'hC52D7374696520766F6C7574706174206E697369206174206665;
        inPKT[558]      = 208'hC52E726D656E74756D2E204E756C6C61206D6F6C657374696520;
        inPKT[559]      = 208'hC52F6E6973692073656420747572706973206D6F6C6573746965;
        inPKT[560]      = 208'hC5302C206E6F6E20696163756C6973206E756E63206661756369;
        inPKT[561]      = 208'hC5316275732E2041656E65616E20696E74657264756D20706861;
        inPKT[562]      = 208'hC532726574726120636F6E73656374657475722E20457469616D;
        inPKT[563]      = 208'hC533206578206F7263692C20696163756C6973206E6F6E206575;
        inPKT[564]      = 208'hC53469736D6F642069642C20756C6C616D636F72706572207363;
        inPKT[565]      = 208'hC535656C65726973717565206F64696F2E0D0A0D0A4E616D2075;
        inPKT[566]      = 208'hC5366C74726963657320656C656966656E64206469616D2C2065;
        inPKT[567]      = 208'hC53767657420736F64616C65732073656D206D61747469732061;
        inPKT[568]      = 208'hC538632E2055742076656E656E61746973206E69626820657520;
        inPKT[569]      = 208'hC5396C65637475732074696E636964756E742064696374756D2E;
        inPKT[570]      = 208'hC53A20566976616D757320637572737573206175677565207175;
        inPKT[571]      = 208'hC53B6973206C6F626F7274697320657569736D6F642E204E756E;
        inPKT[572]      = 208'hC53C6320616C697175616D206469616D20617420616E74652066;
        inPKT[573]      = 208'hC53D6163696C69736973206D6178696D75732E20457469616D20;
        inPKT[574]      = 208'hC53E736564206C6F72656D206D61747469732C20636F6E76616C;
        inPKT[575]      = 208'hC53F6C69732075726E612076697461652C2074656D7075732073;
        inPKT[576]      = 208'hC540656D2E20566976616D7573206567657374617320766F6C75;
        inPKT[577]      = 208'hC541747061742065726F7320657520756C7472696365732E2056;
        inPKT[578]      = 208'hC5426573746962756C756D20756C6C616D636F72706572206572;
        inPKT[579]      = 208'hC5436174206E756E632C206E6F6E2068656E647265726974206F;
        inPKT[580]      = 208'hC54464696F2070656C6C656E7465737175652069642E20467573;
        inPKT[581]      = 208'hC54563652075726E6120697073756D2C206C6163696E69612069;
        inPKT[582]      = 208'hC5466E2073757363697069742076656C2C2073656D7065722069;
        inPKT[583]      = 208'hC5476E206F64696F2E2050656C6C656E74657371756520696420;
        inPKT[584]      = 208'hC5486E696268206E6973692E20416C697175616D20706F727461;
        inPKT[585]      = 208'hC549206E69736C20657420657820696163756C69732074726973;
        inPKT[586]      = 208'hC54A74697175652E20457469616D206D61737361206F7263692C;
        inPKT[587]      = 208'hC54B206567657374617320736564206C6F72656D20717569732C;
        inPKT[588]      = 208'hC54C206469676E697373696D2073656D70657220616E74652E20;
        inPKT[589]      = 208'hC54D53757370656E64697373652074696E636964756E74206E69;
        inPKT[590]      = 208'hC54E73692065782C2073656420766F6C75747061742065737420;
        inPKT[591]      = 208'hC54F7661726975732076697461652E0D0A0D0A5365642073656D;
        inPKT[592]      = 208'hC550706572206C6163696E696120646F6C6F722E204E616D2075;
        inPKT[593]      = 208'hC551742076656C697420696E206C6163757320636F6E73656374;
        inPKT[594]      = 208'hC5526574757220636F6E76616C6C69732070656C6C656E746573;
        inPKT[595]      = 208'hC553717565207365642073656D2E2053757370656E6469737365;
        inPKT[596]      = 208'hC55420636F6E64696D656E74756D20612065726F732069642075;
        inPKT[597]      = 208'hC5556C6C616D636F727065722E204D6F726269206C7563747573;
        inPKT[598]      = 208'hC5562075726E612073697420616D657420657569736D6F642069;
        inPKT[599]      = 208'hC5576163756C69732E2050656C6C656E74657371756520666163;
        inPKT[600]      = 208'hC558696C69736973206D617572697320657520656C656D656E74;
        inPKT[601]      = 208'hC559756D207661726975732E204F72636920766172697573206E;
        inPKT[602]      = 208'hC55A61746F7175652070656E617469627573206574206D61676E;
        inPKT[603]      = 208'hC55B6973206469732070617274757269656E74206D6F6E746573;
        inPKT[604]      = 208'hC55C2C206E61736365747572207269646963756C7573206D7573;
        inPKT[605]      = 208'hC55D2E20446F6E6563206469676E697373696D20612069707375;
        inPKT[606]      = 208'hC55E6D20756C747269636965732076656E656E617469732E2056;
        inPKT[607]      = 208'hC55F6976616D7573206E756E632076656C69742C207665686963;
        inPKT[608]      = 208'hC560756C61207669746165206D617373612075742C20636F6E76;
        inPKT[609]      = 208'hC561616C6C697320636F6E736563746574757220746F72746F72;
        inPKT[610]      = 208'hC5622E205175697371756520616C697175616D2C206E69736C20;
        inPKT[611]      = 208'hC563636F6E67756520626C616E64697420756C74726963696573;
        inPKT[612]      = 208'hC5642C2075726E6120747572706973206D6174746973206D6167;
        inPKT[613]      = 208'hC5656E612C206E6F6E206665726D656E74756D20647569207665;
        inPKT[614]      = 208'hC5666C6974206575207175616D2E0D0A0D0A496E207068617265;
        inPKT[615]      = 208'hC5677472612076656C697420646F6C6F722C2076697461652063;
        inPKT[616]      = 208'hC5687572737573206F7263692066696E696275732074696E6369;
        inPKT[617]      = 208'hC56964756E742E20566976616D757320696420746F72746F7220;
        inPKT[618]      = 208'hC56A72686F6E6375732C207361676974746973206469616D2065;
        inPKT[619]      = 208'hC56B6765742C207072657469756D206D61757269732E20506861;
        inPKT[620]      = 208'hC56C73656C6C757320656C656D656E74756D20656E696D206665;
        inPKT[621]      = 208'hC56D6C69732E204D6175726973206575206E6571756520656765;
        inPKT[622]      = 208'hC56E742070757275732068656E64726572697420677261766964;
        inPKT[623]      = 208'hC56F612E20416C697175616D206C696265726F206E6962682C20;
        inPKT[624]      = 208'hC570636F6E76616C6C69732061206E69736C2065742C2068656E;
        inPKT[625]      = 208'hC57164726572697420766573746962756C756D2066656C69732E;
        inPKT[626]      = 208'hC57220446F6E656320657569736D6F64206665726D656E74756D;
        inPKT[627]      = 208'hC5732074757270697320657520617563746F722E2041656E6561;
        inPKT[628]      = 208'hC5746E20626962656E64756D2074757270697320696E206F6469;
        inPKT[629]      = 208'hC5756F20636F6E76616C6C69732C207669746165207661726975;
        inPKT[630]      = 208'hC57673206578206C616F726565742E2046757363652076656C20;
        inPKT[631]      = 208'hC5776D6920766974616520646F6C6F7220666575676961742076;
        inPKT[632]      = 208'hC578756C707574617465206E6563207574206E756E632E204372;
        inPKT[633]      = 208'hC579617320646170696275732C20616E74652069642076656869;
        inPKT[634]      = 208'hC57A63756C6120616C697175616D2C20656C69742065726F7320;
        inPKT[635]      = 208'hC57B7361676974746973206D692C206E6F6E20656C656966656E;
        inPKT[636]      = 208'hC57C64206578206E756C6C6120656765742076656C69742E2053;
        inPKT[637]      = 208'hC57D757370656E6469737365206964206469616D206475692E20;
        inPKT[638]      = 208'hC57E53757370656E6469737365207072657469756D206A757374;
        inPKT[639]      = 208'hC57F6F20736564206E69626820706F72747469746F722C207665;
        inPKT[640]      = 208'hC5806C20696E74657264756D206D6175726973206D6178696D75;
        inPKT[641]      = 208'hC581732E20557420616C697175616D206C616375732070757275;
        inPKT[642]      = 208'hC582732C2073697420616D657420696D70657264696574206E69;
        inPKT[643]      = 208'hC583626820666575676961742069642E20496E7465676572206C;
        inPKT[644]      = 208'hC5846F72656D206D61757269732C207072657469756D206E6F6E;
        inPKT[645]      = 208'hC585206E6973692065742C20646170696275732066696E696275;
        inPKT[646]      = 208'hC58673206F7263692E0D0A0D0A566573746962756C756D206961;
        inPKT[647]      = 208'hC58763756C69732C206D61676E61206174206D6174746973206D;
        inPKT[648]      = 208'hC5886178696D75732C2061726375206572617420646170696275;
        inPKT[649]      = 208'hC58973206E756E632C206120766172697573206D657475732066;
        inPKT[650]      = 208'hC58A656C697320736564206F7263692E204E756C6C616D206D69;
        inPKT[651]      = 208'hC58B206E6962682C20656C656966656E64206E656320756C7472;
        inPKT[652]      = 208'hC58C69636573206E65632C20636F6E7365637465747572206163;
        inPKT[653]      = 208'hC58D20656E696D2E20536564206C75637475732073656D207175;
        inPKT[654]      = 208'hC58E69732074656D706F7220636F6E6775652E2053757370656E;
        inPKT[655]      = 208'hC58F646973736520706F74656E74692E20457469616D20656765;
        inPKT[656]      = 208'hC59074206C696265726F2076656C69742E204475697320766573;
        inPKT[657]      = 208'hC591746962756C756D20636F6E73657175617420706F7274612E;
        inPKT[658]      = 208'hC592204D617572697320706F72747469746F7220747572706973;
        inPKT[659]      = 208'hC59320696E206D6173736120616C697175616D20636F6E677565;
        inPKT[660]      = 208'hC5942E204E756C6C6120636F6E73656374657475722075726E61;
        inPKT[661]      = 208'hC595206D657475732C20696420696163756C6973206E756E6320;
        inPKT[662]      = 208'hC596756C7472696369657320656765742E204375726162697475;
        inPKT[663]      = 208'hC59772206D6175726973206E657175652C20626962656E64756D;
        inPKT[664]      = 208'hC598207365642065726F732061742C206D6178696D757320756C;
        inPKT[665]      = 208'hC599747269636573207475727069732E0D0A496E74657264756D;
        inPKT[666]      = 208'hC59A206574206D616C6573756164612066616D65732061632061;
        inPKT[667]      = 208'hC59B6E746520697073756D207072696D697320696E2066617563;
        inPKT[668]      = 208'hC59C696275732E2050656C6C656E74657371756520736F6C6C69;
        inPKT[669]      = 208'hC59D6369747564696E20626C616E646974206665726D656E7475;
        inPKT[670]      = 208'hC59E6D2E2050656C6C656E746573717565206E6F6E206C696775;
        inPKT[671]      = 208'hC59F6C6120657520657261742076656E656E6174697320657569;
        inPKT[672]      = 208'hC5A0736D6F642E2050656C6C656E74657371756520736F64616C;
        inPKT[673]      = 208'hC5A1657320766573746962756C756D20636F6E76616C6C69732E;
        inPKT[674]      = 208'hC5A22050726F696E206D6F6C6573746965207072657469756D20;
        inPKT[675]      = 208'hC5A365726F732076656C20656765737461732E204D6F72626920;
        inPKT[676]      = 208'hC5A4736F6C6C696369747564696E207075727573206163206665;
        inPKT[677]      = 208'hC5A5726D656E74756D206D61747469732E204E756E632076656C;
        inPKT[678]      = 208'hC5A62074696E636964756E74206C696265726F2E204E756C6C61;
        inPKT[679]      = 208'hC5A720616C697175657420697073756D206E6563207175616D20;
        inPKT[680]      = 208'hC5A8696D7065726469657420696E74657264756D2E2050726165;
        inPKT[681]      = 208'hC5A973656E74206C6967756C612066656C69732C20696163756C;
        inPKT[682]      = 208'hC5AA697320617420616C69717565742061742C20736167697474;
        inPKT[683]      = 208'hC5AB6973207175697320656C69742E0D0A517569737175652076;
        inPKT[684]      = 208'hC5AC656C20696D70657264696574206E6962682E205068617365;
        inPKT[685]      = 208'hC5AD6C6C75732072757472756D206469676E697373696D207269;
        inPKT[686]      = 208'hC5AE737573206E6F6E2074696E636964756E742E205665737469;
        inPKT[687]      = 208'hC5AF62756C756D206E756E6320697073756D2C2076656E656E61;
        inPKT[688]      = 208'hC5B0746973206567657420706F72746120696E2C20636F6E7365;
        inPKT[689]      = 208'hC5B163746574757220657520657261742E20446F6E6563207665;
        inPKT[690]      = 208'hC5B2686963756C6120616E74652076656C2072686F6E63757320;
        inPKT[691]      = 208'hC5B366617563696275732E2050656C6C656E746573717565206A;
        inPKT[692]      = 208'hC5B47573746F20746F72746F722C20766F6C757470617420696E;
        inPKT[693]      = 208'hC5B5206D61757269732061742C20766172697573207068617265;
        inPKT[694]      = 208'hC5B67472612072697375732E2051756973717565207574206469;
        inPKT[695]      = 208'hC5B7616D2073757363697069742C20736F6C6C69636974756469;
        inPKT[696]      = 208'hC5B86E2073617069656E2065742C20696E74657264756D206C61;
        inPKT[697]      = 208'hC5B96375732E204D6F7262692072697375732073656D2C207065;
        inPKT[698]      = 208'hC5BA6C6C656E7465737175652065742074757270697320696E2C;
        inPKT[699]      = 208'hC5BB20626C616E64697420736F6C6C696369747564696E207365;
        inPKT[700]      = 208'hC5BC6D2E2053656420656666696369747572206C696265726F20;
        inPKT[701]      = 208'hC5BD71756973207072657469756D207072657469756D2E204E75;
        inPKT[702]      = 208'hC5BE6C6C616D20617563746F72207361676974746973206C6F72;
        inPKT[703]      = 208'hC5BF656D2C20616320756C7472696365732061726375206D6178;
        inPKT[704]      = 208'hC5C0696D757320656765742E0D0A566573746962756C756D2076;
        inPKT[705]      = 208'hC5C16F6C7574706174206C6967756C6120617563746F72207365;
        inPKT[706]      = 208'hC5C26D20766976657272612C20756C6C616D636F727065722065;
        inPKT[707]      = 208'hC5C37569736D6F64206E6571756520706F72747469746F722E20;
        inPKT[708]      = 208'hC5C453757370656E64697373652076697665727261207363656C;
        inPKT[709]      = 208'hC5C565726973717565206F64696F2072686F6E63757320766F6C;
        inPKT[710]      = 208'hC5C675747061742E20416C697175616D206572617420766F6C75;
        inPKT[711]      = 208'hC5C7747061742E2053757370656E646973736520706F74656E74;
        inPKT[712]      = 208'hC5C8692E20496E206861632068616269746173736520706C6174;
        inPKT[713]      = 208'hC5C965612064696374756D73742E2050726F696E207574206E75;
        inPKT[714]      = 208'hC5CA6C6C6120757420647569207363656C657269737175652064;
        inPKT[715]      = 208'hC5CB696374756D2E205175697371756520737573636970697420;
        inPKT[716]      = 208'hC5CC6E69626820706F7375657265207175616D2076756C707574;
        inPKT[717]      = 208'hC5CD6174652C206575206C6163696E696120616E746520677261;
        inPKT[718]      = 208'hC5CE766964612E20437572616269747572206D61737361206C6F;
        inPKT[719]      = 208'hC5CF72656D2C206F726E617265206575206D6F6C6C6973206174;
        inPKT[720]      = 208'hC5D02C207068617265747261206E6563206D617373612E204E75;
        inPKT[721]      = 208'hC5D16C6C612066696E6962757320656C656966656E64206F7263;
        inPKT[722]      = 208'hC5D2692073697420616D657420636F6E73656374657475722E20;
        inPKT[723]      = 208'hC5D35365642074656D7075732076697461652061726375206E65;
        inPKT[724]      = 208'hC5D463206665726D656E74756D2E2041656E65616E2070656C6C;
        inPKT[725]      = 208'hC5D5656E74657371756520766974616520646F6C6F7220696E20;
        inPKT[726]      = 208'hC5D6616363756D73616E2E2043726173206469676E697373696D;
        inPKT[727]      = 208'hC5D72076756C707574617465206D6F6C6C69732E204D61757269;
        inPKT[728]      = 208'hC5D87320706F7274612076656E656E617469732072697375732C;
        inPKT[729]      = 208'hC5D92065752074726973746971756520646F6C6F722072757472;
        inPKT[730]      = 208'hC5DA756D20696E2E20467573636520636F6E64696D656E74756D;
        inPKT[731]      = 208'hC5DB206F7263692066656C69732C2073697420616D657420636F;
        inPKT[732]      = 208'hC5DC6E76616C6C6973206C696265726F2074696E636964756E74;
        inPKT[733]      = 208'hC5DD2061632E0D0A566573746962756C756D20696D7065726469;
        inPKT[734]      = 208'hC5DE657420656C69742074656D706F72207175616D2067726176;
        inPKT[735]      = 208'hC5DF6964612C207574206D616C6573756164612074656C6C7573;
        inPKT[736]      = 208'hC5E020696D706572646965742E2050686173656C6C7573206F64;
        inPKT[737]      = 208'hC5E1696F2073656D2C206D61747469732073656420756C747269;
        inPKT[738]      = 208'hC5E26365732061742C20766976657272612076656C206475692E;
        inPKT[739]      = 208'hC5E3204E756E632075726E61206D657475732C206C7563747573;
        inPKT[740]      = 208'hC5E4206163206D6178696D757320696E2C20636F6E7365637465;
        inPKT[741]      = 208'hC5E5747572206E6F6E206E6973692E204E756C6C612073697420;
        inPKT[742]      = 208'hC5E6616D657420626962656E64756D2076656C69742E20446F6E;
        inPKT[743]      = 208'hC5E76563207175697320656E696D206E6F6E2072697375732062;
        inPKT[744]      = 208'hC5E86C616E64697420666163696C697369732071756973206E65;
        inPKT[745]      = 208'hC5E9632072697375732E20437572616269747572206575206573;
        inPKT[746]      = 208'hC5EA74207669746165206C656374757320626C616E6469742061;
        inPKT[747]      = 208'hC5EB6C69717565742E20566573746962756C756D20616E746520;
        inPKT[748]      = 208'hC5EC697073756D207072696D697320696E206661756369627573;
        inPKT[749]      = 208'hC5ED206F726369206C756374757320657420756C747269636573;
        inPKT[750]      = 208'hC5EE20706F737565726520637562696C69612043757261653B20;
        inPKT[751]      = 208'hC5EF566573746962756C756D206163206469676E697373696D20;
        inPKT[752]      = 208'hC5F06E756E632E205175697371756520696E2073616769747469;
        inPKT[753]      = 208'hC5F1732074656C6C75732C2073697420616D6574206665726D65;
        inPKT[754]      = 208'hC5F26E74756D206E6962682E0D0A496E206469676E697373696D;
        inPKT[755]      = 208'hC5F3207269737573207669746165207075727573207665737469;
        inPKT[756]      = 208'hC5F462756C756D2C20617420656C656D656E74756D206E756C6C;
        inPKT[757]      = 208'hC5F56120706F73756572652E20536564206D6174746973206E75;
        inPKT[758]      = 208'hC5F66E63206E6962682E2053757370656E64697373652070656C;
        inPKT[759]      = 208'hC5F76C656E74657371756520706C616365726174207363656C65;
        inPKT[760]      = 208'hC5F87269737175652E2041656E65616E2066657567696174206D;
        inPKT[761]      = 208'hC5F9617572697320696420636F6E677565206C6163696E69612E;
        inPKT[762]      = 208'hC5FA20457469616D207375736369706974206C6967756C612074;
        inPKT[763]      = 208'hC5FB656C6C75732C206120636F6E677565206C65637475732061;
        inPKT[764]      = 208'hC5FC6C697175616D207665686963756C612E2053757370656E64;
        inPKT[765]      = 208'hC5FD69737365206567657420616E74652076656C20656E696D20;
        inPKT[766]      = 208'hC5FE6D616C65737561646120766976657272612E2050726F696E;
        inPKT[767]      = 208'hC5FF2074696E636964756E74206172637520656765742076756C;
        inPKT[768]      = 208'hC50070757461746520616363756D73616E2E20496E2076697461;
        inPKT[769]      = 208'hC50165206469616D206E6962682E204D6F726269206D6178696D;
        inPKT[770]      = 208'hC50275732066656C697320696420636F6E736563746574757220;
        inPKT[771]      = 208'hC503616C697175616D2E204E756C6C6120666163696C6973692E;
        inPKT[772]      = 208'hC5040D0A566573746962756C756D20766573746962756C756D20;
        inPKT[773]      = 208'hC50565666669636974757220746F72746F722073697420616D65;
        inPKT[774]      = 208'hC5067420666163696C697369732E204D616563656E6173206E6F;
        inPKT[775]      = 208'hC5076E2074656C6C7573206F7263692E2050686173656C6C7573;
        inPKT[776]      = 208'hC508206E6F6E206C7563747573206A7573746F2C206174207375;
        inPKT[777]      = 208'hC5097363697069742074656C6C75732E2046757363652068656E;
        inPKT[778]      = 208'hC50A647265726974206E6563206E6962682076656C2063757273;
        inPKT[779]      = 208'hC50B75732E2053757370656E646973736520706F74656E74692E;
        inPKT[780]      = 208'hC50C2044756973206C6967756C612066656C69732C2065666669;
        inPKT[781]      = 208'hC50D63697475722065742076656C69742061742C20666163696C;
        inPKT[782]      = 208'hC50E6973697320636F6E76616C6C6973206A7573746F2E204E75;
        inPKT[783]      = 208'hC50F6C6C616D206C6F626F727469732070656C6C656E74657371;
        inPKT[784]      = 208'hC510756520736F6C6C696369747564696E2E204E616D20736974;
        inPKT[785]      = 208'hC51120616D657420646F6C6F722073697420616D6574206C6563;
        inPKT[786]      = 208'hC51274757320696D7065726469657420636F6E7365717561742E;
        inPKT[787]      = 208'hC51320416C697175616D206C7563747573207363656C65726973;
        inPKT[788]      = 208'hC5147175652070757275732C206964206672696E67696C6C6120;
        inPKT[789]      = 208'hC51573656D20766F6C75747061742061632E205365642074656D;
        inPKT[790]      = 208'hC516706F722C20656E696D206567657420657569736D6F642066;
        inPKT[791]      = 208'hC5176163696C697369732C206E6973692065782073656D706572;
        inPKT[792]      = 208'hC51820697073756D2C20696E207361676974746973206F726369;
        inPKT[793]      = 208'hC519207175616D20696E206C65637475732E2055742076697461;
        inPKT[794]      = 208'hC51A6520656C6974206C6967756C612E204E756E632065676573;
        inPKT[795]      = 208'hC51B7461732C206D6920766974616520696163756C6973206D61;
        inPKT[796]      = 208'hC51C747469732C20647569206E69626820656C656966656E6420;
        inPKT[797]      = 208'hC51D6E69736C2C206567657420706F727461206C696265726F20;
        inPKT[798]      = 208'hC51E6175677565207175697320656E696D2E2053656420736974;
        inPKT[799]      = 208'hC51F20616D65742070756C76696E61722065782C2076656C2070;
        inPKT[800]      = 208'hC520656C6C656E746573717565206C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
