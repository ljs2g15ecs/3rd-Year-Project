//	SIMON_definitions.vh