`include "SIMON_defintions.svh"

module test_SIMON_6496_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 1200
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 144'hE300131211100B0A09080302010000000000;
        inPKT[1]        = 144'hC3014C6F72656D20697073756D20646F6C6F;
        inPKT[2]        = 144'hC302722073697420616D65742C20636F6E73;
        inPKT[3]        = 144'hC30365637465747572206164697069736369;
        inPKT[4]        = 144'hC3046E6720656C69742E2043757261626974;
        inPKT[5]        = 144'hC305757220756C6C616D636F727065722074;
        inPKT[6]        = 144'hC306656D707573206E6973692C2065742070;
        inPKT[7]        = 144'hC3076F73756572652075726E612E2041656E;
        inPKT[8]        = 144'hC30865616E20736564206772617669646120;
        inPKT[9]        = 144'hC3096C616375732E204E756C6C6120666163;
        inPKT[10]       = 144'hC30A696C6973692E204E756C6C612074656D;
        inPKT[11]       = 144'hC30B707573206F726369207175697320656C;
        inPKT[12]       = 144'hC30C697420666575676961742C2076656C20;
        inPKT[13]       = 144'hC30D73656D706572206C656F20696D706572;
        inPKT[14]       = 144'hC30E646965742E204D616563656E61732065;
        inPKT[15]       = 144'hC30F74206E756E6320696E206E6962682066;
        inPKT[16]       = 144'hC3106163696C6973697320636F6E76616C6C;
        inPKT[17]       = 144'hC31169732E2053656420636F6E6775652068;
        inPKT[18]       = 144'hC312656E64726572697420696163756C6973;
        inPKT[19]       = 144'hC3132E20566976616D757320766568696375;
        inPKT[20]       = 144'hC3146C61206C7563747573206573742C2076;
        inPKT[21]       = 144'hC31569746165207375736369706974206E69;
        inPKT[22]       = 144'hC316736C20706F72747469746F722061632E;
        inPKT[23]       = 144'hC3170D0A0D0A446F6E6563206D6F6C657374;
        inPKT[24]       = 144'hC31869652073617069656E2069642076756C;
        inPKT[25]       = 144'hC31970757461746520766573746962756C75;
        inPKT[26]       = 144'hC31A6D2E204E756C6C6120696E206C696775;
        inPKT[27]       = 144'hC31B6C61206672696E67696C6C612C20756C;
        inPKT[28]       = 144'hC31C6C616D636F727065722075726E612065;
        inPKT[29]       = 144'hC31D742C20706F72747469746F72206C6563;
        inPKT[30]       = 144'hC31E7475732E205175697371756520626C61;
        inPKT[31]       = 144'hC31F6E646974206575206D61757269732061;
        inPKT[32]       = 144'hC320632068656E6472657269742E204E756C;
        inPKT[33]       = 144'hC3216C612076656E656E617469732C206D65;
        inPKT[34]       = 144'hC322747573206574206C7563747573206672;
        inPKT[35]       = 144'hC323696E67696C6C612C206E696268207665;
        inPKT[36]       = 144'hC3246C697420756C6C616D636F7270657220;
        inPKT[37]       = 144'hC3256469616D2C2065676574206566666963;
        inPKT[38]       = 144'hC3266974757220697073756D207475727069;
        inPKT[39]       = 144'hC32773206174206E6962682E205574206567;
        inPKT[40]       = 144'hC3286574207072657469756D2065726F732C;
        inPKT[41]       = 144'hC32920656765742064696374756D206C6163;
        inPKT[42]       = 144'hC32A75732E204D616563656E617320757420;
        inPKT[43]       = 144'hC32B656E696D2065782E2041656E65616E20;
        inPKT[44]       = 144'hC32C76697461652073656D7065722066656C;
        inPKT[45]       = 144'hC32D69732C2073656420756C747269636965;
        inPKT[46]       = 144'hC32E732072697375732E20446F6E65632063;
        inPKT[47]       = 144'hC32F6F6E7365637465747572206D69206E69;
        inPKT[48]       = 144'hC330736C2C20617420637572737573206970;
        inPKT[49]       = 144'hC33173756D206772617669646120612E2050;
        inPKT[50]       = 144'hC332686173656C6C75732073697420616D65;
        inPKT[51]       = 144'hC33374206D61676E612076656C2069707375;
        inPKT[52]       = 144'hC3346D206567657374617320706F7274612E;
        inPKT[53]       = 144'hC33520566976616D7573206C756374757320;
        inPKT[54]       = 144'hC336656E696D20656765742074656D706F72;
        inPKT[55]       = 144'hC3372073616769747469732E20416C697175;
        inPKT[56]       = 144'hC338616D20626962656E64756D2073656D20;
        inPKT[57]       = 144'hC3396120636F6E7365637465747572206566;
        inPKT[58]       = 144'hC33A666963697475722E20446F6E65632073;
        inPKT[59]       = 144'hC33B63656C6572697371756520616C697175;
        inPKT[60]       = 144'hC33C616D206375727375732E204375726162;
        inPKT[61]       = 144'hC33D697475722073697420616D6574206269;
        inPKT[62]       = 144'hC33E62656E64756D20656C69742E20536564;
        inPKT[63]       = 144'hC33F206469616D206A7573746F2C20696163;
        inPKT[64]       = 144'hC340756C69732071756973206E756C6C6120;
        inPKT[65]       = 144'hC34176697461652C20616C697175616D2065;
        inPKT[66]       = 144'hC3427569736D6F642066656C69732E0D0A0D;
        inPKT[67]       = 144'hC3430A50726F696E20646170696275732C20;
        inPKT[68]       = 144'hC3446469616D2076756C7075746174652066;
        inPKT[69]       = 144'hC34572696E67696C6C61206D616C65737561;
        inPKT[70]       = 144'hC34664612C206A7573746F20707572757320;
        inPKT[71]       = 144'hC347636F6D6D6F646F20646F6C6F722C2075;
        inPKT[72]       = 144'hC348742064696374756D2065726174206E75;
        inPKT[73]       = 144'hC3496E632072757472756D2075726E612E20;
        inPKT[74]       = 144'hC34A4E756C6C612067726176696461207572;
        inPKT[75]       = 144'hC34B6E6120766974616520696D7065726469;
        inPKT[76]       = 144'hC34C6574206C616F726565742E2050656C6C;
        inPKT[77]       = 144'hC34D656E7465737175652072686F6E637573;
        inPKT[78]       = 144'hC34E20626962656E64756D206E6962682C20;
        inPKT[79]       = 144'hC34F6964206D6F6C6C6973206469616D2073;
        inPKT[80]       = 144'hC350757363697069742061632E2050656C6C;
        inPKT[81]       = 144'hC351656E7465737175652076656C20696163;
        inPKT[82]       = 144'hC352756C6973206475692E204D6F72626920;
        inPKT[83]       = 144'hC353617420616C6971756574206D61737361;
        inPKT[84]       = 144'hC3542E2050726F696E207669746165206F72;
        inPKT[85]       = 144'hC3556E617265206F64696F2C206575207675;
        inPKT[86]       = 144'hC3566C70757461746520697073756D2E2050;
        inPKT[87]       = 144'hC357726F696E206C6F626F727469732C2073;
        inPKT[88]       = 144'hC358656D206E656320657569736D6F642074;
        inPKT[89]       = 144'hC359696E636964756E742C20617567756520;
        inPKT[90]       = 144'hC35A6D6175726973207363656C6572697371;
        inPKT[91]       = 144'hC35B7565206D61676E612C20657420706F73;
        inPKT[92]       = 144'hC35C75657265206D69206E69736C206E6563;
        inPKT[93]       = 144'hC35D206E6973692E20467573636520656C69;
        inPKT[94]       = 144'hC35E74206E657175652C2076617269757320;
        inPKT[95]       = 144'hC35F6574206672696E67696C6C6120766974;
        inPKT[96]       = 144'hC36061652C207661726975732076656C206E;
        inPKT[97]       = 144'hC361657175652E204E756C6C612065742074;
        inPKT[98]       = 144'hC362656D707573206A7573746F2E204D6F72;
        inPKT[99]       = 144'hC363626920756C6C616D636F727065722073;
        inPKT[100]      = 144'hC3647573636970697420636F6E6775652E20;
        inPKT[101]      = 144'hC36553656420656C656966656E64206F6469;
        inPKT[102]      = 144'hC3666F206163207375736369706974206469;
        inPKT[103]      = 144'hC367676E697373696D2E2051756973717565;
        inPKT[104]      = 144'hC36820616E746520656E696D2C20626C616E;
        inPKT[105]      = 144'hC36964697420696E20636F6E736571756174;
        inPKT[106]      = 144'hC36A2061632C20696E74657264756D207669;
        inPKT[107]      = 144'hC36B7461652070757275732E204D61757269;
        inPKT[108]      = 144'hC36C7320657569736D6F6420706F73756572;
        inPKT[109]      = 144'hC36D65206C65637475732E20566976616D75;
        inPKT[110]      = 144'hC36E7320696E74657264756D207175616D20;
        inPKT[111]      = 144'hC36F65752073656D70657220666175636962;
        inPKT[112]      = 144'hC37075732E0D0A0D0A496E206D6F6C657374;
        inPKT[113]      = 144'hC3716965206E756C6C6120616E74652C2061;
        inPKT[114]      = 144'hC3726320696E74657264756D206D61676E61;
        inPKT[115]      = 144'hC37320636F6E64696D656E74756D20636F6E;
        inPKT[116]      = 144'hC37464696D656E74756D2E20447569732075;
        inPKT[117]      = 144'hC3756C7472696369657320736F64616C6573;
        inPKT[118]      = 144'hC376206E756C6C612C2073697420616D6574;
        inPKT[119]      = 144'hC37720756C6C616D636F72706572206F6469;
        inPKT[120]      = 144'hC3786F207072657469756D206E65632E2046;
        inPKT[121]      = 144'hC37975736365207365642072697375732070;
        inPKT[122]      = 144'hC37A656C6C656E7465737175652C20636F6E;
        inPKT[123]      = 144'hC37B76616C6C69732073656D20656765742C;
        inPKT[124]      = 144'hC37C2068656E64726572697420657261742E;
        inPKT[125]      = 144'hC37D204D6F72626920736F64616C65732076;
        inPKT[126]      = 144'hC37E65686963756C61206C6F626F72746973;
        inPKT[127]      = 144'hC37F2E2041656E65616E206120746F72746F;
        inPKT[128]      = 144'hC38072206375727375732C207363656C6572;
        inPKT[129]      = 144'hC3816973717565206C6967756C6120706F72;
        inPKT[130]      = 144'hC382747469746F722C206567657374617320;
        inPKT[131]      = 144'hC38365726F732E20447569732074696E6369;
        inPKT[132]      = 144'hC38464756E7420746F72746F722069642070;
        inPKT[133]      = 144'hC3856F737565726520677261766964612E20;
        inPKT[134]      = 144'hC386496E20636F6E76616C6C6973206D6920;
        inPKT[135]      = 144'hC387696420697073756D206D616C65737561;
        inPKT[136]      = 144'hC38864612C2075742064696374756D206572;
        inPKT[137]      = 144'hC3896F7320696D706572646965742E205072;
        inPKT[138]      = 144'hC38A6F696E20756C6C616D636F727065722C;
        inPKT[139]      = 144'hC38B206D6175726973206964207661726975;
        inPKT[140]      = 144'hC38C7320636F6E6775652C2065726F732073;
        inPKT[141]      = 144'hC38D617069656E2072686F6E637573206D69;
        inPKT[142]      = 144'hC38E2C20617420617563746F72206E657175;
        inPKT[143]      = 144'hC38F652061726375206C616F726565742064;
        inPKT[144]      = 144'hC39069616D2E0D0A0D0A467573636520706F;
        inPKT[145]      = 144'hC39172747469746F72206C696265726F2061;
        inPKT[146]      = 144'hC3927263752C206C6163696E69612068656E;
        inPKT[147]      = 144'hC393647265726974206469616D20636F6E76;
        inPKT[148]      = 144'hC394616C6C6973207365642E205068617365;
        inPKT[149]      = 144'hC3956C6C7573206E6F6E2074757270697320;
        inPKT[150]      = 144'hC39670686172657472612C20756C6C616D63;
        inPKT[151]      = 144'hC3976F72706572206E657175652076656C2C;
        inPKT[152]      = 144'hC39820736F6C6C696369747564696E207665;
        inPKT[153]      = 144'hC3996C69742E2050656C6C656E7465737175;
        inPKT[154]      = 144'hC39A65206861626974616E74206D6F726269;
        inPKT[155]      = 144'hC39B207472697374697175652073656E6563;
        inPKT[156]      = 144'hC39C747573206574206E6574757320657420;
        inPKT[157]      = 144'hC39D6D616C6573756164612066616D657320;
        inPKT[158]      = 144'hC39E61632074757270697320656765737461;
        inPKT[159]      = 144'hC39F732E204E616D206E6563207361706965;
        inPKT[160]      = 144'hC3A06E206D6F6C65737469652C2064696374;
        inPKT[161]      = 144'hC3A1756D206D6173736120656765742C2065;
        inPKT[162]      = 144'hC3A2676573746173206F64696F2E20457469;
        inPKT[163]      = 144'hC3A3616D20617263752073617069656E2C20;
        inPKT[164]      = 144'hC3A47072657469756D2061206D6F6C6C6973;
        inPKT[165]      = 144'hC3A520612C2076756C707574617465206E6F;
        inPKT[166]      = 144'hC3A66E20657261742E205574207669746165;
        inPKT[167]      = 144'hC3A7206E696268206C6F626F72746973206C;
        inPKT[168]      = 144'hC3A865637475732066617563696275732070;
        inPKT[169]      = 144'hC3A96F7274612065752073697420616D6574;
        inPKT[170]      = 144'hC3AA206E69736C2E204D6F72626920706F72;
        inPKT[171]      = 144'hC3AB747469746F722076656C697420657520;
        inPKT[172]      = 144'hC3AC646F6C6F72206C616F726565742C2073;
        inPKT[173]      = 144'hC3AD697420616D657420696D706572646965;
        inPKT[174]      = 144'hC3AE7420656E696D20736F64616C65732E20;
        inPKT[175]      = 144'hC3AF4E756C6C616D20756C6C616D636F7270;
        inPKT[176]      = 144'hC3B06572207475727069732061742070656C;
        inPKT[177]      = 144'hC3B16C656E74657371756520766172697573;
        inPKT[178]      = 144'hC3B22E20566976616D757320657520696D70;
        inPKT[179]      = 144'hC3B3657264696574206E657175652E205365;
        inPKT[180]      = 144'hC3B464207175697320617563746F7220616E;
        inPKT[181]      = 144'hC3B574652E204D61757269732073656D7065;
        inPKT[182]      = 144'hC3B67220697073756D207365642064756920;
        inPKT[183]      = 144'hC3B7706F73756572652C20617420616C6971;
        inPKT[184]      = 144'hC3B875616D206D6574757320656C65696665;
        inPKT[185]      = 144'hC3B96E642E204E756C6C616D207472697374;
        inPKT[186]      = 144'hC3BA6971756520656C656966656E64206572;
        inPKT[187]      = 144'hC3BB6F732C2065676574206665726D656E74;
        inPKT[188]      = 144'hC3BC756D20697073756D20656C656D656E74;
        inPKT[189]      = 144'hC3BD756D206E65632E0D0A0D0A50656C6C65;
        inPKT[190]      = 144'hC3BE6E7465737175652068656E6472657269;
        inPKT[191]      = 144'hC3BF7420626962656E64756D206C6967756C;
        inPKT[192]      = 144'hC3C0612C20657420736F64616C6573206D61;
        inPKT[193]      = 144'hC3C1676E61206461706962757320696E2E20;
        inPKT[194]      = 144'hC3C2496E20616C697175657420746F72746F;
        inPKT[195]      = 144'hC3C372206567657420636F6E736563746574;
        inPKT[196]      = 144'hC3C4757220636F6E73656374657475722E20;
        inPKT[197]      = 144'hC3C551756973717565207472697374697175;
        inPKT[198]      = 144'hC3C66520726973757320657261742C206574;
        inPKT[199]      = 144'hC3C720616C697175657420656C697420616C;
        inPKT[200]      = 144'hC3C869717565742065752E20496E74656765;
        inPKT[201]      = 144'hC3C972206E6F6E206D61676E6120696E2066;
        inPKT[202]      = 144'hC3CA656C697320706F72747469746F722073;
        inPKT[203]      = 144'hC3CB616769747469732E2051756973717565;
        inPKT[204]      = 144'hC3CC2076697665727261206F726369206163;
        inPKT[205]      = 144'hC3CD2072757472756D206C616F726565742E;
        inPKT[206]      = 144'hC3CE2041656E65616E20636F6E76616C6C69;
        inPKT[207]      = 144'hC3CF732064696374756D207475727069732C;
        inPKT[208]      = 144'hC3D02065742066696E696275732073617069;
        inPKT[209]      = 144'hC3D1656E20636F6E67756520696E2E205365;
        inPKT[210]      = 144'hC3D26420612065726174206F726E6172652C;
        inPKT[211]      = 144'hC3D3206D6F6C6C6973206E69736C2061632C;
        inPKT[212]      = 144'hC3D4206469676E697373696D206E65717565;
        inPKT[213]      = 144'hC3D52E2051756973717565206D616C657375;
        inPKT[214]      = 144'hC3D661646120706F73756572652074757270;
        inPKT[215]      = 144'hC3D7697320657520756C6C616D636F727065;
        inPKT[216]      = 144'hC3D8722E20446F6E65632076697665727261;
        inPKT[217]      = 144'hC3D920626962656E64756D206E756E632C20;
        inPKT[218]      = 144'hC3DA64696374756D20696D70657264696574;
        inPKT[219]      = 144'hC3DB206E65717565206D6178696D75732069;
        inPKT[220]      = 144'hC3DC6E2E20446F6E656320757420756C7472;
        inPKT[221]      = 144'hC3DD6963657320646F6C6F722E2056697661;
        inPKT[222]      = 144'hC3DE6D757320736564206175677565207072;
        inPKT[223]      = 144'hC3DF657469756D2C20766F6C757470617420;
        inPKT[224]      = 144'hC3E0657261742061632C20706F7274612064;
        inPKT[225]      = 144'hC3E169616D2E204D617572697320696E2070;
        inPKT[226]      = 144'hC3E27572757320756C747269636965732C20;
        inPKT[227]      = 144'hC3E37375736369706974206469616D207365;
        inPKT[228]      = 144'hC3E4642C2074696E636964756E7420656E69;
        inPKT[229]      = 144'hC3E56D2E20446F6E6563207175697320706F;
        inPKT[230]      = 144'hC3E67375657265206E6962682E20496E2068;
        inPKT[231]      = 144'hC3E761632068616269746173736520706C61;
        inPKT[232]      = 144'hC3E87465612064696374756D73742E0D0A0D;
        inPKT[233]      = 144'hC3E90A4D6F726269206F726E617265206A75;
        inPKT[234]      = 144'hC3EA73746F206174207175616D2066617563;
        inPKT[235]      = 144'hC3EB696275732C2073697420616D6574206D;
        inPKT[236]      = 144'hC3EC6F6C6573746965206C656F2063757273;
        inPKT[237]      = 144'hC3ED75732E204D6175726973206C616F7265;
        inPKT[238]      = 144'hC3EE657420616E74652061206D6574757320;
        inPKT[239]      = 144'hC3EF65666669636974757220766172697573;
        inPKT[240]      = 144'hC3F02E205365642076656C206F7263692073;
        inPKT[241]      = 144'hC3F161676974746973206E756E6320626C61;
        inPKT[242]      = 144'hC3F26E64697420636F6E7365717561742E20;
        inPKT[243]      = 144'hC3F35072616573656E74206D616C65737561;
        inPKT[244]      = 144'hC3F46461206E657175652071756973206469;
        inPKT[245]      = 144'hC3F56374756D206469676E697373696D2E20;
        inPKT[246]      = 144'hC3F6446F6E656320666163696C6973697320;
        inPKT[247]      = 144'hC3F773697420616D65742076656C69742065;
        inPKT[248]      = 144'hC3F875206C6F626F727469732E204E756C6C;
        inPKT[249]      = 144'hC3F9616D20626C616E64697420656C656D65;
        inPKT[250]      = 144'hC3FA6E74756D206D61757269732C20766974;
        inPKT[251]      = 144'hC3FB616520656C656D656E74756D20646F6C;
        inPKT[252]      = 144'hC3FC6F722068656E64726572697420766974;
        inPKT[253]      = 144'hC3FD61652E204675736365206D6F6C657374;
        inPKT[254]      = 144'hC3FE69652C20656C697420757420616C6971;
        inPKT[255]      = 144'hC3FF75657420766F6C75747061742C206E65;
        inPKT[256]      = 144'hC3007175652076656C697420707265746975;
        inPKT[257]      = 144'hC3016D2061756775652C206672696E67696C;
        inPKT[258]      = 144'hC3026C6120636F6E64696D656E74756D206A;
        inPKT[259]      = 144'hC3037573746F2073617069656E2061206A75;
        inPKT[260]      = 144'hC30473746F2E2050686173656C6C75732071;
        inPKT[261]      = 144'hC30575697320617563746F72206C6F72656D;
        inPKT[262]      = 144'hC3062C20696E20616C697175616D206E756E;
        inPKT[263]      = 144'hC307632E20557420656C656966656E642061;
        inPKT[264]      = 144'hC3086E7465206574206E697369206D6F6C65;
        inPKT[265]      = 144'hC3097374696520636F6E76616C6C69732069;
        inPKT[266]      = 144'hC30A642065742073656D2E20536564206163;
        inPKT[267]      = 144'hC30B20626962656E64756D20617263752E20;
        inPKT[268]      = 144'hC30C467573636520766573746962756C756D;
        inPKT[269]      = 144'hC30D206E756E6320656765742074656C6C75;
        inPKT[270]      = 144'hC30E73206665726D656E74756D2C206E6563;
        inPKT[271]      = 144'hC30F2072686F6E637573206D617373612063;
        inPKT[272]      = 144'hC3106F6D6D6F646F2E204D616563656E6173;
        inPKT[273]      = 144'hC311206964206E756E63206E6F6E20657820;
        inPKT[274]      = 144'hC312766573746962756C756D206F726E6172;
        inPKT[275]      = 144'hC31365207574206E65632065726F732E2041;
        inPKT[276]      = 144'hC3146C697175616D20656666696369747572;
        inPKT[277]      = 144'hC31520636F6D6D6F646F206469616D206964;
        inPKT[278]      = 144'hC316206C6F626F727469732E205365642061;
        inPKT[279]      = 144'hC317632074656D706F72206C65637475732E;
        inPKT[280]      = 144'hC318204E756E6320656C656D656E74756D20;
        inPKT[281]      = 144'hC3197574206C65637475732061632074696E;
        inPKT[282]      = 144'hC31A636964756E742E20557420696163756C;
        inPKT[283]      = 144'hC31B6973206E756C6C612071756973206578;
        inPKT[284]      = 144'hC31C20656C656D656E74756D2C20616C6971;
        inPKT[285]      = 144'hC31D7565742073656D706572206D61676E61;
        inPKT[286]      = 144'hC31E20656C656966656E642E0D0A0D0A4375;
        inPKT[287]      = 144'hC31F7261626974757220746F72746F72206E;
        inPKT[288]      = 144'hC32069736C2C20756C747269636965732069;
        inPKT[289]      = 144'hC3216E206E657175652061632C2061636375;
        inPKT[290]      = 144'hC3226D73616E20636F6E736571756174206D;
        inPKT[291]      = 144'hC323657475732E204D616563656E6173206D;
        inPKT[292]      = 144'hC324617373612073617069656E2C206D6174;
        inPKT[293]      = 144'hC32574697320696E2076656E656E61746973;
        inPKT[294]      = 144'hC3262073697420616D65742C20617563746F;
        inPKT[295]      = 144'hC327722073697420616D657420656E696D2E;
        inPKT[296]      = 144'hC328204E756E63207669746165206D657475;
        inPKT[297]      = 144'hC3297320636F6D6D6F646F2C206D61747469;
        inPKT[298]      = 144'hC32A73206D617373612073697420616D6574;
        inPKT[299]      = 144'hC32B2C20766172697573206C6F72656D2E20;
        inPKT[300]      = 144'hC32C4E756E6320696E20656C697420656C69;
        inPKT[301]      = 144'hC32D742E204E756E63206F726E6172652063;
        inPKT[302]      = 144'hC32E6F6E7365637465747572206D61676E61;
        inPKT[303]      = 144'hC32F2C2073697420616D657420706F727474;
        inPKT[304]      = 144'hC33069746F7220617263752072686F6E6375;
        inPKT[305]      = 144'hC331732065752E2053757370656E64697373;
        inPKT[306]      = 144'hC33265207363656C6572697371756520756C;
        inPKT[307]      = 144'hC33374726963696573206578206120616C69;
        inPKT[308]      = 144'hC3347175616D2E2053757370656E64697373;
        inPKT[309]      = 144'hC335652072757472756D20736F6C6C696369;
        inPKT[310]      = 144'hC336747564696E206E756E632C206E6F6E20;
        inPKT[311]      = 144'hC337636F6E76616C6C697320747572706973;
        inPKT[312]      = 144'hC338206C616F726565742073697420616D65;
        inPKT[313]      = 144'hC339742E2041656E65616E20612066696E69;
        inPKT[314]      = 144'hC33A627573206D61757269732C2071756973;
        inPKT[315]      = 144'hC33B20637572737573206E756E632E20496E;
        inPKT[316]      = 144'hC33C2066657567696174206475692076656C;
        inPKT[317]      = 144'hC33D2075726E612073656D70657220666175;
        inPKT[318]      = 144'hC33E63696275732E204D617572697320756C;
        inPKT[319]      = 144'hC33F74726963696573206174207475727069;
        inPKT[320]      = 144'hC3407320656765742070656C6C656E746573;
        inPKT[321]      = 144'hC3417175652E205072616573656E74207369;
        inPKT[322]      = 144'hC3427420616D6574206C6967756C6120636F;
        inPKT[323]      = 144'hC3436E76616C6C69732C20656C656D656E74;
        inPKT[324]      = 144'hC344756D206E756C6C6120756C6C616D636F;
        inPKT[325]      = 144'hC345727065722C20616C697175616D207572;
        inPKT[326]      = 144'hC3466E612E20457469616D207175616D2065;
        inPKT[327]      = 144'hC3476C69742C20706F737565726520757420;
        inPKT[328]      = 144'hC3487175616D20656765742C2066696E6962;
        inPKT[329]      = 144'hC349757320736F6C6C696369747564696E20;
        inPKT[330]      = 144'hC34A6E756C6C612E20496E20737573636970;
        inPKT[331]      = 144'hC34B697420656E696D2065742065726F7320;
        inPKT[332]      = 144'hC34C66696E696275732C207574207363656C;
        inPKT[333]      = 144'hC34D657269737175652074656C6C75732066;
        inPKT[334]      = 144'hC34E6575676961742E204375726162697475;
        inPKT[335]      = 144'hC34F72206E6F6E206D617373612076617269;
        inPKT[336]      = 144'hC350757320646F6C6F722067726176696461;
        inPKT[337]      = 144'hC35120656C656D656E74756D207175697320;
        inPKT[338]      = 144'hC35275742066656C69732E2050686173656C;
        inPKT[339]      = 144'hC3536C757320657569736D6F642069707375;
        inPKT[340]      = 144'hC3546D20656765742076656C6974206C6F62;
        inPKT[341]      = 144'hC3556F727469732C206567657420706F7274;
        inPKT[342]      = 144'hC35661206D61757269732074656D7075732E;
        inPKT[343]      = 144'hC3572053656420696D706572646965742076;
        inPKT[344]      = 144'hC3586F6C75747061742074656C6C75732065;
        inPKT[345]      = 144'hC359752074696E636964756E742E0D0A0D0A;
        inPKT[346]      = 144'hC35A55742076656C206D69206174206D6574;
        inPKT[347]      = 144'hC35B7573206672696E67696C6C6120677261;
        inPKT[348]      = 144'hC35C766964612E205072616573656E742065;
        inPKT[349]      = 144'hC35D726F73206E6962682C20637572737573;
        inPKT[350]      = 144'hC35E20656765737461732074696E63696475;
        inPKT[351]      = 144'hC35F6E7420736F64616C65732C207363656C;
        inPKT[352]      = 144'hC36065726973717565206E65632066656C69;
        inPKT[353]      = 144'hC361732E20496E746567657220696D706572;
        inPKT[354]      = 144'hC36264696574206D616C657375616461206E;
        inPKT[355]      = 144'hC36369736C20616C69717565742076656E65;
        inPKT[356]      = 144'hC3646E617469732E20496E74656765722073;
        inPKT[357]      = 144'hC365656420706F72747469746F7220697073;
        inPKT[358]      = 144'hC366756D2E20496E746567657220636F6D6D;
        inPKT[359]      = 144'hC3676F646F206665756769617420746F7274;
        inPKT[360]      = 144'hC3686F722C206575206C6F626F7274697320;
        inPKT[361]      = 144'hC369617567756520656C656D656E74756D20;
        inPKT[362]      = 144'hC36A73697420616D65742E20446F6E656320;
        inPKT[363]      = 144'hC36B766573746962756C756D206C6967756C;
        inPKT[364]      = 144'hC36C612061756775652C2065742066696E69;
        inPKT[365]      = 144'hC36D627573206172637520706F7274612069;
        inPKT[366]      = 144'hC36E6E2E204E756C6C612073656D2074656C;
        inPKT[367]      = 144'hC36F6C75732C20756C6C616D636F72706572;
        inPKT[368]      = 144'hC3702061742063757273757320612C20706F;
        inPKT[369]      = 144'hC3717274612073697420616D6574206D6167;
        inPKT[370]      = 144'hC3726E612E204E756E632076697461652069;
        inPKT[371]      = 144'hC3736D706572646965742070757275732C20;
        inPKT[372]      = 144'hC3746E656320736F6C6C696369747564696E;
        inPKT[373]      = 144'hC3752074656C6C75732E20416C697175616D;
        inPKT[374]      = 144'hC376206572617420766F6C75747061742E20;
        inPKT[375]      = 144'hC377536564206964206D61676E6120636F6D;
        inPKT[376]      = 144'hC3786D6F646F2C206C75637475732076656C;
        inPKT[377]      = 144'hC379697420717569732C20657569736D6F64;
        inPKT[378]      = 144'hC37A20656E696D2E20496E7465676572206D;
        inPKT[379]      = 144'hC37B617474697320736F64616C6573206665;
        inPKT[380]      = 144'hC37C726D656E74756D2E2051756973717565;
        inPKT[381]      = 144'hC37D20736564206672696E67696C6C61206C;
        inPKT[382]      = 144'hC37E6F72656D2E2043726173207665686963;
        inPKT[383]      = 144'hC37F756C612074656D707573207361706965;
        inPKT[384]      = 144'hC3806E20757420636F6E6775652E20447569;
        inPKT[385]      = 144'hC381732073617069656E20656E696D2C2070;
        inPKT[386]      = 144'hC3826F727461206E6563206C656F2069642C;
        inPKT[387]      = 144'hC3832065666669636974757220706F737565;
        inPKT[388]      = 144'hC3847265206C696265726F2E204E756C6C61;
        inPKT[389]      = 144'hC3856D2061632074656D706F72206D657475;
        inPKT[390]      = 144'hC386732E205365642076656C207475727069;
        inPKT[391]      = 144'hC3877320666575676961742C20696163756C;
        inPKT[392]      = 144'hC388697320617567756520717569732C2074;
        inPKT[393]      = 144'hC389696E636964756E74207475727069732E;
        inPKT[394]      = 144'hC38A0D0A0D0A566976616D757320706F7375;
        inPKT[395]      = 144'hC38B65726520706F72747469746F72206175;
        inPKT[396]      = 144'hC38C6775652C207661726975732061636375;
        inPKT[397]      = 144'hC38D6D73616E20656C69742076756C707574;
        inPKT[398]      = 144'hC38E61746520656765742E20517569737175;
        inPKT[399]      = 144'hC38F6520736564206D616C65737561646120;
        inPKT[400]      = 144'hC3906E69736C2E20496E74657264756D2065;
        inPKT[401]      = 144'hC39174206D616C6573756164612066616D65;
        inPKT[402]      = 144'hC3927320616320616E746520697073756D20;
        inPKT[403]      = 144'hC3937072696D697320696E20666175636962;
        inPKT[404]      = 144'hC39475732E204E756E632074757270697320;
        inPKT[405]      = 144'hC3956469616D2C2073757363697069742061;
        inPKT[406]      = 144'hC396632065726F732076656C2C2074656D70;
        inPKT[407]      = 144'hC39775732076656E656E6174697320697073;
        inPKT[408]      = 144'hC398756D2E2044756973206C756374757320;
        inPKT[409]      = 144'hC39972686F6E637573206D617373612E2046;
        inPKT[410]      = 144'hC39A75736365207574206C6163696E696120;
        inPKT[411]      = 144'hC39B7475727069732E20566976616D757320;
        inPKT[412]      = 144'hC39C72757472756D2074656C6C7573206175;
        inPKT[413]      = 144'hC39D6775652C206174206F726E617265206E;
        inPKT[414]      = 144'hC39E69736C20666163696C69736973206574;
        inPKT[415]      = 144'hC39F2E204E756E6320736564206E69736920;
        inPKT[416]      = 144'hC3A072697375732E20496E74656765722065;
        inPKT[417]      = 144'hC3A16C656D656E74756D206D617572697320;
        inPKT[418]      = 144'hC3A27175616D2C207574207665686963756C;
        inPKT[419]      = 144'hC3A361206D617572697320636F6E67756520;
        inPKT[420]      = 144'hC3A465752E0D0A0D0A467573636520612074;
        inPKT[421]      = 144'hC3A5656C6C75732073697420616D65742065;
        inPKT[422]      = 144'hC3A6726174206665726D656E74756D207363;
        inPKT[423]      = 144'hC3A7656C657269737175652E204375726162;
        inPKT[424]      = 144'hC3A86974757220696E2076656C6974206174;
        inPKT[425]      = 144'hC3A920656E696D206C6163696E6961207665;
        inPKT[426]      = 144'hC3AA686963756C61206163206964206A7573;
        inPKT[427]      = 144'hC3AB746F2E2050726F696E206E6F6E20646F;
        inPKT[428]      = 144'hC3AC6C6F72206566666963697475722C2074;
        inPKT[429]      = 144'hC3AD696E636964756E74206F64696F206575;
        inPKT[430]      = 144'hC3AE2C20666175636962757320656E696D2E;
        inPKT[431]      = 144'hC3AF2050656C6C656E746573717565206461;
        inPKT[432]      = 144'hC3B07069627573206F726369206163206C6F;
        inPKT[433]      = 144'hC3B172656D20696163756C69732C20736974;
        inPKT[434]      = 144'hC3B220616D657420626C616E646974206172;
        inPKT[435]      = 144'hC3B36375207472697374697175652E204165;
        inPKT[436]      = 144'hC3B46E65616E207472697374697175652074;
        inPKT[437]      = 144'hC3B56F72746F72206E6563206A7573746F20;
        inPKT[438]      = 144'hC3B6616C697175616D2C20696E2070726574;
        inPKT[439]      = 144'hC3B769756D2066656C6973206D6F6C657374;
        inPKT[440]      = 144'hC3B869652E205365642065742074656D7075;
        inPKT[441]      = 144'hC3B9732061756775652E204E756C6C612066;
        inPKT[442]      = 144'hC3BA72696E67696C6C6120656C656966656E;
        inPKT[443]      = 144'hC3BB6420697073756D207669766572726120;
        inPKT[444]      = 144'hC3BC6375727375732E20416C697175616D20;
        inPKT[445]      = 144'hC3BD6D6178696D7573206665726D656E7475;
        inPKT[446]      = 144'hC3BE6D206E69626820616320616363756D73;
        inPKT[447]      = 144'hC3BF616E2E204E756C6C6120666163696C69;
        inPKT[448]      = 144'hC3C073692E20566573746962756C756D2066;
        inPKT[449]      = 144'hC3C16163696C69736973206C656F20656765;
        inPKT[450]      = 144'hC3C2737461732073656D206D617474697320;
        inPKT[451]      = 144'hC3C3636F6E6775652E204D61757269732076;
        inPKT[452]      = 144'hC3C469746165206578206174207269737573;
        inPKT[453]      = 144'hC3C5206461706962757320656C656966656E;
        inPKT[454]      = 144'hC3C6642E20496E7465676572207574206572;
        inPKT[455]      = 144'hC3C76F7320636F6E6775652C20706F727474;
        inPKT[456]      = 144'hC3C869746F7220616E7465206E6F6E2C2069;
        inPKT[457]      = 144'hC3C96E74657264756D20646F6C6F722E0D0A;
        inPKT[458]      = 144'hC3CA0D0A566573746962756C756D20656C65;
        inPKT[459]      = 144'hC3CB6966656E64206D617572697320657520;
        inPKT[460]      = 144'hC3CC6E6973692064696374756D2067726176;
        inPKT[461]      = 144'hC3CD6964612E2044756973206D6F6C6C6973;
        inPKT[462]      = 144'hC3CE206469616D2076656C20656E696D2074;
        inPKT[463]      = 144'hC3CF656D7075732C20766974616520646170;
        inPKT[464]      = 144'hC3D069627573206D61737361207361676974;
        inPKT[465]      = 144'hC3D17469732E204E756C6C61207574206175;
        inPKT[466]      = 144'hC3D263746F7220746F72746F722E204D6F72;
        inPKT[467]      = 144'hC3D3626920736564206C6F72656D2075726E;
        inPKT[468]      = 144'hC3D4612E204675736365206D61747469732C;
        inPKT[469]      = 144'hC3D5206D61676E6120616320636F6E64696D;
        inPKT[470]      = 144'hC3D6656E74756D20666575676961742C206D;
        inPKT[471]      = 144'hC3D76173736120647569206D6178696D7573;
        inPKT[472]      = 144'hC3D8206E756C6C612C20657520616C697175;
        inPKT[473]      = 144'hC3D96574206E65717565206D617572697320;
        inPKT[474]      = 144'hC3DA6120657261742E205175697371756520;
        inPKT[475]      = 144'hC3DB617563746F722065737420757420696E;
        inPKT[476]      = 144'hC3DC74657264756D20636F6E736563746574;
        inPKT[477]      = 144'hC3DD75722E20446F6E656320656765742064;
        inPKT[478]      = 144'hC3DE69676E697373696D20746F72746F722C;
        inPKT[479]      = 144'hC3DF2068656E647265726974206D61747469;
        inPKT[480]      = 144'hC3E07320657261742E2050656C6C656E7465;
        inPKT[481]      = 144'hC3E173717565206861626974616E74206D6F;
        inPKT[482]      = 144'hC3E272626920747269737469717565207365;
        inPKT[483]      = 144'hC3E36E6563747573206574206E6574757320;
        inPKT[484]      = 144'hC3E46574206D616C6573756164612066616D;
        inPKT[485]      = 144'hC3E565732061632074757270697320656765;
        inPKT[486]      = 144'hC3E6737461732E2051756973717565206F72;
        inPKT[487]      = 144'hC3E76E617265207661726975732074656D70;
        inPKT[488]      = 144'hC3E875732E0D0A0D0A4D6F72626920727574;
        inPKT[489]      = 144'hC3E972756D20616E7465206E6962682C2061;
        inPKT[490]      = 144'hC3EA2076697665727261206E756C6C612068;
        inPKT[491]      = 144'hC3EB656E64726572697420696E2E2050726F;
        inPKT[492]      = 144'hC3EC696E2073757363697069742065676573;
        inPKT[493]      = 144'hC3ED74617320657261742C20757420617563;
        inPKT[494]      = 144'hC3EE746F72206F726369206D617474697320;
        inPKT[495]      = 144'hC3EF612E2050656C6C656E74657371756520;
        inPKT[496]      = 144'hC3F06C7563747573206672696E67696C6C61;
        inPKT[497]      = 144'hC3F120656C6974207574206C6163696E6961;
        inPKT[498]      = 144'hC3F22E205574206574206D61737361206E75;
        inPKT[499]      = 144'hC3F36C6C612E20536564206174206672696E;
        inPKT[500]      = 144'hC3F467696C6C61206C6F72656D2E2050726F;
        inPKT[501]      = 144'hC3F5696E206772617669646120616363756D;
        inPKT[502]      = 144'hC3F673616E20726973757320736564206269;
        inPKT[503]      = 144'hC3F762656E64756D2E204D616563656E6173;
        inPKT[504]      = 144'hC3F8206D616C657375616461206F64696F20;
        inPKT[505]      = 144'hC3F975742076656C697420657569736D6F64;
        inPKT[506]      = 144'hC3FA20646170696275732E0D0A0D0A457469;
        inPKT[507]      = 144'hC3FB616D20636F6E677565206D6174746973;
        inPKT[508]      = 144'hC3FC20696163756C69732E204D6175726973;
        inPKT[509]      = 144'hC3FD20766974616520656666696369747572;
        inPKT[510]      = 144'hC3FE2073656D2E205365642070756C76696E;
        inPKT[511]      = 144'hC3FF617220646F6C6F72207574206D692065;
        inPKT[512]      = 144'hC3007569736D6F642068656E647265726974;
        inPKT[513]      = 144'hC3012E204E756C6C616D2061742067726176;
        inPKT[514]      = 144'hC30269646120646F6C6F722E204D6F726269;
        inPKT[515]      = 144'hC303206C656F207475727069732C20636F6E;
        inPKT[516]      = 144'hC304677565206E656320616C697175616D20;
        inPKT[517]      = 144'hC30575742C20636F6D6D6F646F20696E206E;
        inPKT[518]      = 144'hC306756E632E204E756C6C61206174206661;
        inPKT[519]      = 144'hC307756369627573206C656F2C2065752066;
        inPKT[520]      = 144'hC308657567696174206C616375732E204675;
        inPKT[521]      = 144'hC309736365206E6F6E206567657374617320;
        inPKT[522]      = 144'hC30A7475727069732E205175697371756520;
        inPKT[523]      = 144'hC30B766974616520697073756D206D692E20;
        inPKT[524]      = 144'hC30C4E756E63206E6F6E206F726369207369;
        inPKT[525]      = 144'hC30D7420616D6574206E6973692076617269;
        inPKT[526]      = 144'hC30E757320706F72747469746F7220696E20;
        inPKT[527]      = 144'hC30F76756C70757461746520746F72746F72;
        inPKT[528]      = 144'hC3102E204E756E6320636F6E76616C6C6973;
        inPKT[529]      = 144'hC3112067726176696461206469616D206120;
        inPKT[530]      = 144'hC312756C747269636965732E205175697371;
        inPKT[531]      = 144'hC3137565206575206A7573746F20636F6E64;
        inPKT[532]      = 144'hC314696D656E74756D2C2076617269757320;
        inPKT[533]      = 144'hC3156469616D2076656C2C20766573746962;
        inPKT[534]      = 144'hC316756C756D206D617373612E0D0A0D0A50;
        inPKT[535]      = 144'hC317656C6C656E7465737175652070656C6C;
        inPKT[536]      = 144'hC318656E7465737175652073617069656E20;
        inPKT[537]      = 144'hC3196E657175652C20617563746F72206D61;
        inPKT[538]      = 144'hC31A6C65737561646120657261742068656E;
        inPKT[539]      = 144'hC31B647265726974206E65632E204E756C6C;
        inPKT[540]      = 144'hC31C6120706C616365726174206469616D20;
        inPKT[541]      = 144'hC31D68656E647265726974206D6173736120;
        inPKT[542]      = 144'hC31E626962656E64756D2C2061206D6F6C65;
        inPKT[543]      = 144'hC31F737469652066656C69732068656E6472;
        inPKT[544]      = 144'hC320657269742E204D617572697320657569;
        inPKT[545]      = 144'hC321736D6F642076656E656E61746973206A;
        inPKT[546]      = 144'hC3227573746F2C20757420617563746F7220;
        inPKT[547]      = 144'hC323656C697420616C69717565742075742E;
        inPKT[548]      = 144'hC32420467573636520616C69717565742C20;
        inPKT[549]      = 144'hC3257175616D207574206469676E69737369;
        inPKT[550]      = 144'hC3266D2068656E6472657269742C206D6175;
        inPKT[551]      = 144'hC32772697320747572706973206469676E69;
        inPKT[552]      = 144'hC3287373696D20746F72746F722C20656765;
        inPKT[553]      = 144'hC329742070656C6C656E7465737175652076;
        inPKT[554]      = 144'hC32A656C6974206F726369206E6563207175;
        inPKT[555]      = 144'hC32B616D2E204E756E632065676573746173;
        inPKT[556]      = 144'hC32C2070656C6C656E746573717565207269;
        inPKT[557]      = 144'hC32D7375732E204375726162697475722073;
        inPKT[558]      = 144'hC32E757363697069742074656D707573206C;
        inPKT[559]      = 144'hC32F616375732C2065676574207072657469;
        inPKT[560]      = 144'hC330756D20656C69742074696E636964756E;
        inPKT[561]      = 144'hC33174206E6F6E2E20437261732075726E61;
        inPKT[562]      = 144'hC332206C6F72656D2C20706C616365726174;
        inPKT[563]      = 144'hC33320766F6C757470617420696D70657264;
        inPKT[564]      = 144'hC3346965742073697420616D65742C206567;
        inPKT[565]      = 144'hC33565737461732076656C206F7263692E0D;
        inPKT[566]      = 144'hC3360A0D0A50656C6C656E74657371756520;
        inPKT[567]      = 144'hC337736F64616C6573206665726D656E7475;
        inPKT[568]      = 144'hC3386D206E69736C2C206174206672696E67;
        inPKT[569]      = 144'hC339696C6C61206475692073656D70657220;
        inPKT[570]      = 144'hC33A6665726D656E74756D2E204E756C6C61;
        inPKT[571]      = 144'hC33B6D20706C6163657261742076656C206D;
        inPKT[572]      = 144'hC33C692068656E64726572697420656C656D;
        inPKT[573]      = 144'hC33D656E74756D2E20457469616D206E6F6E;
        inPKT[574]      = 144'hC33E20697073756D2065782E204E616D2061;
        inPKT[575]      = 144'hC33F63207363656C65726973717565206E69;
        inPKT[576]      = 144'hC34062682C2076656C20666163696C697369;
        inPKT[577]      = 144'hC34173206D692E20446F6E65632065676573;
        inPKT[578]      = 144'hC342746173206C616F726565742065726F73;
        inPKT[579]      = 144'hC3432C206567657420766F6C757470617420;
        inPKT[580]      = 144'hC3446D657475732E205072616573656E7420;
        inPKT[581]      = 144'hC345616363756D73616E20626962656E6475;
        inPKT[582]      = 144'hC3466D206E69736C206E65632076656E656E;
        inPKT[583]      = 144'hC347617469732E205365642072757472756D;
        inPKT[584]      = 144'hC348206D6920612073757363697069742070;
        inPKT[585]      = 144'hC349686172657472612E2053656420736974;
        inPKT[586]      = 144'hC34A20616D657420696E74657264756D2074;
        inPKT[587]      = 144'hC34B75727069732E20416C697175616D2065;
        inPKT[588]      = 144'hC34C75206E69626820746F72746F722E2044;
        inPKT[589]      = 144'hC34D6F6E6563206661756369627573206461;
        inPKT[590]      = 144'hC34E7069627573206E6973692C2073656420;
        inPKT[591]      = 144'hC34F6C616F72656574206F72636920736365;
        inPKT[592]      = 144'hC3506C6572697371756520696E2E0D0A0D0A;
        inPKT[593]      = 144'hC3514D617572697320696E2066656C697320;
        inPKT[594]      = 144'hC3526665726D656E74756D2C20636F6E7661;
        inPKT[595]      = 144'hC3536C6C69732061756775652076656C2C20;
        inPKT[596]      = 144'hC354706F7375657265206D692E2050656C6C;
        inPKT[597]      = 144'hC355656E746573717565207363656C657269;
        inPKT[598]      = 144'hC356737175652072686F6E637573206A7573;
        inPKT[599]      = 144'hC357746F2C2065752070756C76696E617220;
        inPKT[600]      = 144'hC358656E696D2070756C76696E6172207665;
        inPKT[601]      = 144'hC3596C2E204D616563656E61732070686172;
        inPKT[602]      = 144'hC35A65747261206C696265726F206D61676E;
        inPKT[603]      = 144'hC35B612C20616320736F6C6C696369747564;
        inPKT[604]      = 144'hC35C696E206C656F206D6F6C6C6973206E6F;
        inPKT[605]      = 144'hC35D6E2E204E756C6C6120656C656D656E74;
        inPKT[606]      = 144'hC35E756D206F726E61726520656765737461;
        inPKT[607]      = 144'hC35F732E20436C61737320617074656E7420;
        inPKT[608]      = 144'hC36074616369746920736F63696F73717520;
        inPKT[609]      = 144'hC3616164206C69746F726120746F72717565;
        inPKT[610]      = 144'hC3626E742070657220636F6E75626961206E;
        inPKT[611]      = 144'hC3636F737472612C2070657220696E636570;
        inPKT[612]      = 144'hC364746F732068696D656E61656F732E2050;
        inPKT[613]      = 144'hC36572616573656E74206175677565206D61;
        inPKT[614]      = 144'hC366757269732C2072686F6E637573207175;
        inPKT[615]      = 144'hC367697320657374206E6F6E2C206D6F6C6C;
        inPKT[616]      = 144'hC368697320636F6E76616C6C69732066656C;
        inPKT[617]      = 144'hC36969732E2053757370656E646973736520;
        inPKT[618]      = 144'hC36A666163696C697369732C206F72636920;
        inPKT[619]      = 144'hC36B7669746165206C6163696E6961207465;
        inPKT[620]      = 144'hC36C6D706F722C206C656374757320736170;
        inPKT[621]      = 144'hC36D69656E206D6174746973207269737573;
        inPKT[622]      = 144'hC36E2C206E6F6E2073616769747469732065;
        inPKT[623]      = 144'hC36F6C6974206E657175652071756973206A;
        inPKT[624]      = 144'hC3707573746F2E20446F6E6563206D616C65;
        inPKT[625]      = 144'hC3717375616461206C6163696E6961206475;
        inPKT[626]      = 144'hC372692E2050686173656C6C75732068656E;
        inPKT[627]      = 144'hC373647265726974206D6175726973206D61;
        inPKT[628]      = 144'hC374757269732C20736564206672696E6769;
        inPKT[629]      = 144'hC3756C6C61206C696265726F206672696E67;
        inPKT[630]      = 144'hC376696C6C6120696E2E2053656420617420;
        inPKT[631]      = 144'hC3776C6967756C6120696E206A7573746F20;
        inPKT[632]      = 144'hC37866696E696275732076756C7075746174;
        inPKT[633]      = 144'hC379652E204E756E6320637572737573206E;
        inPKT[634]      = 144'hC37A657175652073697420616D6574206172;
        inPKT[635]      = 144'hC37B63752074696E636964756E742C207669;
        inPKT[636]      = 144'hC37C7461652070686172657472612073656D;
        inPKT[637]      = 144'hC37D20706F72747469746F722E20416C6971;
        inPKT[638]      = 144'hC37E75616D206D61747469732C206A757374;
        inPKT[639]      = 144'hC37F6F206E6F6E20657569736D6F6420636F;
        inPKT[640]      = 144'hC3806E76616C6C69732C206E756E63206D69;
        inPKT[641]      = 144'hC38120636F6E736571756174206573742C20;
        inPKT[642]      = 144'hC3826E656320736F6C6C696369747564696E;
        inPKT[643]      = 144'hC383206C65637475732073617069656E2076;
        inPKT[644]      = 144'hC384656C206F64696F2E20496E2074656D70;
        inPKT[645]      = 144'hC3856F72206572617420646F6C6F722C2073;
        inPKT[646]      = 144'hC3866564207665686963756C612075726E61;
        inPKT[647]      = 144'hC38720636F6E736571756174207365642E0D;
        inPKT[648]      = 144'hC3880A0D0A4E616D2072686F6E6375732069;
        inPKT[649]      = 144'hC38964206D6175726973206E656320646967;
        inPKT[650]      = 144'hC38A6E697373696D2E20496E20696D706572;
        inPKT[651]      = 144'hC38B6469657420756C747269636573206572;
        inPKT[652]      = 144'hC38C6174206E656320736F6C6C6963697475;
        inPKT[653]      = 144'hC38D64696E2E20496E746567657220736564;
        inPKT[654]      = 144'hC38E20636F6E64696D656E74756D2065726F;
        inPKT[655]      = 144'hC38F732E20446F6E65632065676574206E75;
        inPKT[656]      = 144'hC3906E63206964206D617572697320747269;
        inPKT[657]      = 144'hC39173746971756520706F72747469746F72;
        inPKT[658]      = 144'hC392206C616F72656574207669746165206D;
        inPKT[659]      = 144'hC393657475732E204E756C6C612066616369;
        inPKT[660]      = 144'hC3946C6973692E204E756C6C616D20657520;
        inPKT[661]      = 144'hC3956C616375732061206469616D20747269;
        inPKT[662]      = 144'hC3967374697175652065676573746173206E;
        inPKT[663]      = 144'hC3976F6E20696163756C6973206D65747573;
        inPKT[664]      = 144'hC3982E20416C697175616D20696E2074656D;
        inPKT[665]      = 144'hC399706F7220657261742C20696420636F6E;
        inPKT[666]      = 144'hC39A677565206D617373612E20566976616D;
        inPKT[667]      = 144'hC39B75732076656C20746F72746F72207669;
        inPKT[668]      = 144'hC39C746165206E69626820636F6D6D6F646F;
        inPKT[669]      = 144'hC39D206C6F626F7274697320717569732061;
        inPKT[670]      = 144'hC39E20697073756D2E2050726F696E20766F;
        inPKT[671]      = 144'hC39F6C7574706174207175616D206E6F6E20;
        inPKT[672]      = 144'hC3A066656C69732074656D7075732C206964;
        inPKT[673]      = 144'hC3A120706F737565726520646F6C6F722074;
        inPKT[674]      = 144'hC3A2656D706F722E205072616573656E7420;
        inPKT[675]      = 144'hC3A376697461652074696E636964756E7420;
        inPKT[676]      = 144'hC3A473617069656E2E204D616563656E6173;
        inPKT[677]      = 144'hC3A520666163696C69736973206D61747469;
        inPKT[678]      = 144'hC3A67320616E746520717569732076617269;
        inPKT[679]      = 144'hC3A775732E20446F6E65632070656C6C656E;
        inPKT[680]      = 144'hC3A87465737175652065726F732066657567;
        inPKT[681]      = 144'hC3A96961742074696E636964756E7420636F;
        inPKT[682]      = 144'hC3AA6E64696D656E74756D2E2050726F696E;
        inPKT[683]      = 144'hC3AB20666175636962757320766F6C757470;
        inPKT[684]      = 144'hC3AC6174206D692073656420736167697474;
        inPKT[685]      = 144'hC3AD69732E0D0A0D0A447569732067726176;
        inPKT[686]      = 144'hC3AE69646120656C656D656E74756D20696E;
        inPKT[687]      = 144'hC3AF74657264756D2E2050726F696E207369;
        inPKT[688]      = 144'hC3B07420616D6574207175616D206C696775;
        inPKT[689]      = 144'hC3B16C612E2050686173656C6C757320636F;
        inPKT[690]      = 144'hC3B26D6D6F646F2C2075726E6120696E2063;
        inPKT[691]      = 144'hC3B36F6E67756520766F6C75747061742C20;
        inPKT[692]      = 144'hC3B46C6967756C6120657820706861726574;
        inPKT[693]      = 144'hC3B57261206C6967756C612C20696E206469;
        inPKT[694]      = 144'hC3B66374756D206D61676E61206F72636920;
        inPKT[695]      = 144'hC3B76E6563206D61757269732E204E756E63;
        inPKT[696]      = 144'hC3B820617563746F7220636F6E7365637465;
        inPKT[697]      = 144'hC3B974757220766F6C75747061742E204D6F;
        inPKT[698]      = 144'hC3BA7262692074696E636964756E74206E69;
        inPKT[699]      = 144'hC3BB626820757420656E696D206566666963;
        inPKT[700]      = 144'hC3BC6974757220677261766964612E204375;
        inPKT[701]      = 144'hC3BD72616269747572207669746165207175;
        inPKT[702]      = 144'hC3BE616D2065726F732E2044756973206672;
        inPKT[703]      = 144'hC3BF696E67696C6C6120616320746F72746F;
        inPKT[704]      = 144'hC3C07220696E2074696E636964756E742E20;
        inPKT[705]      = 144'hC3C14E756E632076656C206D617572697320;
        inPKT[706]      = 144'hC3C272697375732E20446F6E656320656C65;
        inPKT[707]      = 144'hC3C36966656E64206C6967756C6120736167;
        inPKT[708]      = 144'hC3C46974746973206E6973692066696E6962;
        inPKT[709]      = 144'hC3C575732C2061207363656C657269737175;
        inPKT[710]      = 144'hC3C665206C696265726F2070656C6C656E74;
        inPKT[711]      = 144'hC3C765737175652E20566573746962756C75;
        inPKT[712]      = 144'hC3C86D20747269737469717565206D617373;
        inPKT[713]      = 144'hC3C961206E6962682C206174207665737469;
        inPKT[714]      = 144'hC3CA62756C756D206D61676E612066696E69;
        inPKT[715]      = 144'hC3CB6275732065752E0D0A0D0A4375726162;
        inPKT[716]      = 144'hC3CC6974757220696D706572646965742070;
        inPKT[717]      = 144'hC3CD757275732065676574206E756E632075;
        inPKT[718]      = 144'hC3CE6C7472696365732C2076697461652076;
        inPKT[719]      = 144'hC3CF656E656E61746973206D617373612063;
        inPKT[720]      = 144'hC3D06F6D6D6F646F2E2050656C6C656E7465;
        inPKT[721]      = 144'hC3D173717565206861626974616E74206D6F;
        inPKT[722]      = 144'hC3D272626920747269737469717565207365;
        inPKT[723]      = 144'hC3D36E6563747573206574206E6574757320;
        inPKT[724]      = 144'hC3D46574206D616C6573756164612066616D;
        inPKT[725]      = 144'hC3D565732061632074757270697320656765;
        inPKT[726]      = 144'hC3D6737461732E20496E206665726D656E74;
        inPKT[727]      = 144'hC3D7756D2061742075726E61206E6F6E2063;
        inPKT[728]      = 144'hC3D86F6E76616C6C69732E20446F6E656320;
        inPKT[729]      = 144'hC3D96163206175677565206A7573746F2E20;
        inPKT[730]      = 144'hC3DA496E20617420656C6974206574206172;
        inPKT[731]      = 144'hC3DB6375206D6178696D7573206C75637475;
        inPKT[732]      = 144'hC3DC732E20467573636520657569736D6F64;
        inPKT[733]      = 144'hC3DD206E756E63206E65632076656E656E61;
        inPKT[734]      = 144'hC3DE74697320617563746F722E204C6F7265;
        inPKT[735]      = 144'hC3DF6D20697073756D20646F6C6F72207369;
        inPKT[736]      = 144'hC3E07420616D65742C20636F6E7365637465;
        inPKT[737]      = 144'hC3E17475722061646970697363696E672065;
        inPKT[738]      = 144'hC3E26C69742E20446F6E6563206469637475;
        inPKT[739]      = 144'hC3E36D2074656D706F722072757472756D2E;
        inPKT[740]      = 144'hC3E42053656420656C656966656E64206469;
        inPKT[741]      = 144'hC3E5616D206964206D6173736120696D7065;
        inPKT[742]      = 144'hC3E672646965742C206163206F726E617265;
        inPKT[743]      = 144'hC3E7206C696265726F20656C656966656E64;
        inPKT[744]      = 144'hC3E82E204D616563656E6173206F726E6172;
        inPKT[745]      = 144'hC3E965206D65747573206E756C6C612C2073;
        inPKT[746]      = 144'hC3EA697420616D6574206665726D656E7475;
        inPKT[747]      = 144'hC3EB6D20656C697420616C697175616D2069;
        inPKT[748]      = 144'hC3EC642E20446F6E656320756C7472696365;
        inPKT[749]      = 144'hC3ED7320746F72746F7220617420616E7465;
        inPKT[750]      = 144'hC3EE2068656E6472657269742C2065752073;
        inPKT[751]      = 144'hC3EF61676974746973206A7573746F20756C;
        inPKT[752]      = 144'hC3F07472696365732E0D0A0D0A5072616573;
        inPKT[753]      = 144'hC3F1656E74206C7563747573207072657469;
        inPKT[754]      = 144'hC3F2756D206E657175652C2073697420616D;
        inPKT[755]      = 144'hC3F365742070656C6C656E74657371756520;
        inPKT[756]      = 144'hC3F46D617572697320656C656D656E74756D;
        inPKT[757]      = 144'hC3F5206E6F6E2E20557420626C616E646974;
        inPKT[758]      = 144'hC3F6207068617265747261206F64696F206E;
        inPKT[759]      = 144'hC3F76F6E20657569736D6F642E2051756973;
        inPKT[760]      = 144'hC3F8717565207669746165206C656F20616C;
        inPKT[761]      = 144'hC3F9697175616D2C20736F64616C65732074;
        inPKT[762]      = 144'hC3FA656C6C75732069642C20696163756C69;
        inPKT[763]      = 144'hC3FB73206D61757269732E204E616D206566;
        inPKT[764]      = 144'hC3FC6669636974757220696E207075727573;
        inPKT[765]      = 144'hC3FD2073656420616363756D73616E2E204D;
        inPKT[766]      = 144'hC3FE616563656E61732073697420616D6574;
        inPKT[767]      = 144'hC3FF206375727375732066656C69732E2051;
        inPKT[768]      = 144'hC3007569737175652066617563696275732C;
        inPKT[769]      = 144'hC3012064756920657420617563746F72206C;
        inPKT[770]      = 144'hC30275637475732C20616E74652065726174;
        inPKT[771]      = 144'hC30320706F73756572652065726F732C2075;
        inPKT[772]      = 144'hC3047420636F6E76616C6C6973206D657475;
        inPKT[773]      = 144'hC30573206C6563747573207669746165206C;
        inPKT[774]      = 144'hC306656F2E2053757370656E646973736520;
        inPKT[775]      = 144'hC307706F74656E74692E2043726173206574;
        inPKT[776]      = 144'hC30820646F6C6F72206E6F6E2075726E6120;
        inPKT[777]      = 144'hC3097363656C657269737175652074726973;
        inPKT[778]      = 144'hC30A74697175652E20437261732072757472;
        inPKT[779]      = 144'hC30B756D206E65632076656C697420616320;
        inPKT[780]      = 144'hC30C73616769747469732E20446F6E656320;
        inPKT[781]      = 144'hC30D656C656966656E642C206C6163757320;
        inPKT[782]      = 144'hC30E7365642067726176696461206D616C65;
        inPKT[783]      = 144'hC30F73756164612C20657820616E74652070;
        inPKT[784]      = 144'hC3106C616365726174206C65637475732C20;
        inPKT[785]      = 144'hC3116567657420636F6E677565206D617373;
        inPKT[786]      = 144'hC31261206D65747573206964206C61637573;
        inPKT[787]      = 144'hC3132E2053757370656E6469737365206964;
        inPKT[788]      = 144'hC3142072757472756D206C65637475732E20;
        inPKT[789]      = 144'hC3154675736365206D6178696D7573207365;
        inPKT[790]      = 144'hC31664206C6967756C612073656420766976;
        inPKT[791]      = 144'hC317657272612E204E616D206C7563747573;
        inPKT[792]      = 144'hC318206469616D20616E74652C2076697461;
        inPKT[793]      = 144'hC31965206F726E617265206E657175652076;
        inPKT[794]      = 144'hC31A617269757320656765742E0D0A0D0A50;
        inPKT[795]      = 144'hC31B656C6C656E7465737175652061742065;
        inPKT[796]      = 144'hC31C6C6974206E6962682E20566573746962;
        inPKT[797]      = 144'hC31D756C756D20616E746520697073756D20;
        inPKT[798]      = 144'hC31E7072696D697320696E20666175636962;
        inPKT[799]      = 144'hC31F7573206F726369206C75637475732065;
        inPKT[800]      = 144'hC3207420756C74726963657320706F737565;
        inPKT[801]      = 144'hC321726520637562696C6961204375726165;
        inPKT[802]      = 144'hC3223B204375726162697475722066617563;
        inPKT[803]      = 144'hC32369627573206469616D206C656F2C206E;
        inPKT[804]      = 144'hC324656320657569736D6F642073656D2065;
        inPKT[805]      = 144'hC32566666963697475722075742E20557420;
        inPKT[806]      = 144'hC3267665686963756C612061756775652061;
        inPKT[807]      = 144'hC32763206C696265726F20696163756C6973;
        inPKT[808]      = 144'hC3282C206E656320656C656966656E642065;
        inPKT[809]      = 144'hC3297820706F7274612E204D6F7262692068;
        inPKT[810]      = 144'hC32A656E6472657269742067726176696461;
        inPKT[811]      = 144'hC32B2074696E636964756E742E2050726165;
        inPKT[812]      = 144'hC32C73656E7420646F6C6F72206C61637573;
        inPKT[813]      = 144'hC32D2C2074656D707573206575206672696E;
        inPKT[814]      = 144'hC32E67696C6C612073697420616D65742C20;
        inPKT[815]      = 144'hC32F656C656966656E6420696E206E756C6C;
        inPKT[816]      = 144'hC330612E204E756C6C61206D6F6C6C697320;
        inPKT[817]      = 144'hC33165676574206D61676E61206E65632068;
        inPKT[818]      = 144'hC332656E6472657269742E20416C69717561;
        inPKT[819]      = 144'hC3336D20636F6E76616C6C69732073656D20;
        inPKT[820]      = 144'hC33476697461652073617069656E20646963;
        inPKT[821]      = 144'hC33574756D2C20757420766573746962756C;
        inPKT[822]      = 144'hC336756D206C6F72656D206672696E67696C;
        inPKT[823]      = 144'hC3376C612E20446F6E65632074656C6C7573;
        inPKT[824]      = 144'hC338206C696265726F2C2066657567696174;
        inPKT[825]      = 144'hC3392075742066696E69627573206E65632C;
        inPKT[826]      = 144'hC33A20616C697175616D2073697420616D65;
        inPKT[827]      = 144'hC33B74206F7263692E204E756E6320737573;
        inPKT[828]      = 144'hC33C6369706974206E69736C206574206F72;
        inPKT[829]      = 144'hC33D6E61726520766573746962756C756D2E;
        inPKT[830]      = 144'hC33E204E756C6C616D206C6F626F72746973;
        inPKT[831]      = 144'hC33F2073617069656E206A7573746F2C2073;
        inPKT[832]      = 144'hC340697420616D6574206469676E69737369;
        inPKT[833]      = 144'hC3416D206E756C6C6120636F6E64696D656E;
        inPKT[834]      = 144'hC34274756D20696E2E20536564206D6F6C65;
        inPKT[835]      = 144'hC3437374696520766F6C7574706174206E69;
        inPKT[836]      = 144'hC3447369206174206665726D656E74756D2E;
        inPKT[837]      = 144'hC345204E756C6C61206D6F6C657374696520;
        inPKT[838]      = 144'hC3466E697369207365642074757270697320;
        inPKT[839]      = 144'hC3476D6F6C65737469652C206E6F6E206961;
        inPKT[840]      = 144'hC34863756C6973206E756E63206661756369;
        inPKT[841]      = 144'hC3496275732E2041656E65616E20696E7465;
        inPKT[842]      = 144'hC34A7264756D20706861726574726120636F;
        inPKT[843]      = 144'hC34B6E73656374657475722E20457469616D;
        inPKT[844]      = 144'hC34C206578206F7263692C20696163756C69;
        inPKT[845]      = 144'hC34D73206E6F6E20657569736D6F64206964;
        inPKT[846]      = 144'hC34E2C20756C6C616D636F72706572207363;
        inPKT[847]      = 144'hC34F656C65726973717565206F64696F2E0D;
        inPKT[848]      = 144'hC3500A0D0A4E616D20756C74726963657320;
        inPKT[849]      = 144'hC351656C656966656E64206469616D2C2065;
        inPKT[850]      = 144'hC35267657420736F64616C65732073656D20;
        inPKT[851]      = 144'hC3536D61747469732061632E205574207665;
        inPKT[852]      = 144'hC3546E656E61746973206E69626820657520;
        inPKT[853]      = 144'hC3556C65637475732074696E636964756E74;
        inPKT[854]      = 144'hC3562064696374756D2E20566976616D7573;
        inPKT[855]      = 144'hC35720637572737573206175677565207175;
        inPKT[856]      = 144'hC3586973206C6F626F727469732065756973;
        inPKT[857]      = 144'hC3596D6F642E204E756E6320616C69717561;
        inPKT[858]      = 144'hC35A6D206469616D20617420616E74652066;
        inPKT[859]      = 144'hC35B6163696C69736973206D6178696D7573;
        inPKT[860]      = 144'hC35C2E20457469616D20736564206C6F7265;
        inPKT[861]      = 144'hC35D6D206D61747469732C20636F6E76616C;
        inPKT[862]      = 144'hC35E6C69732075726E612076697461652C20;
        inPKT[863]      = 144'hC35F74656D7075732073656D2E2056697661;
        inPKT[864]      = 144'hC3606D7573206567657374617320766F6C75;
        inPKT[865]      = 144'hC361747061742065726F7320657520756C74;
        inPKT[866]      = 144'hC36272696365732E20566573746962756C75;
        inPKT[867]      = 144'hC3636D20756C6C616D636F72706572206572;
        inPKT[868]      = 144'hC3646174206E756E632C206E6F6E2068656E;
        inPKT[869]      = 144'hC365647265726974206F64696F2070656C6C;
        inPKT[870]      = 144'hC366656E7465737175652069642E20467573;
        inPKT[871]      = 144'hC36763652075726E6120697073756D2C206C;
        inPKT[872]      = 144'hC3686163696E696120696E20737573636970;
        inPKT[873]      = 144'hC36969742076656C2C2073656D7065722069;
        inPKT[874]      = 144'hC36A6E206F64696F2E2050656C6C656E7465;
        inPKT[875]      = 144'hC36B73717565206964206E696268206E6973;
        inPKT[876]      = 144'hC36C692E20416C697175616D20706F727461;
        inPKT[877]      = 144'hC36D206E69736C2065742065782069616375;
        inPKT[878]      = 144'hC36E6C6973207472697374697175652E2045;
        inPKT[879]      = 144'hC36F7469616D206D61737361206F7263692C;
        inPKT[880]      = 144'hC370206567657374617320736564206C6F72;
        inPKT[881]      = 144'hC371656D20717569732C206469676E697373;
        inPKT[882]      = 144'hC372696D2073656D70657220616E74652E20;
        inPKT[883]      = 144'hC37353757370656E64697373652074696E63;
        inPKT[884]      = 144'hC3746964756E74206E6973692065782C2073;
        inPKT[885]      = 144'hC375656420766F6C75747061742065737420;
        inPKT[886]      = 144'hC3767661726975732076697461652E0D0A0D;
        inPKT[887]      = 144'hC3770A5365642073656D706572206C616369;
        inPKT[888]      = 144'hC3786E696120646F6C6F722E204E616D2075;
        inPKT[889]      = 144'hC379742076656C697420696E206C61637573;
        inPKT[890]      = 144'hC37A20636F6E736563746574757220636F6E;
        inPKT[891]      = 144'hC37B76616C6C69732070656C6C656E746573;
        inPKT[892]      = 144'hC37C717565207365642073656D2E20537573;
        inPKT[893]      = 144'hC37D70656E646973736520636F6E64696D65;
        inPKT[894]      = 144'hC37E6E74756D20612065726F732069642075;
        inPKT[895]      = 144'hC37F6C6C616D636F727065722E204D6F7262;
        inPKT[896]      = 144'hC38069206C75637475732075726E61207369;
        inPKT[897]      = 144'hC3817420616D657420657569736D6F642069;
        inPKT[898]      = 144'hC3826163756C69732E2050656C6C656E7465;
        inPKT[899]      = 144'hC3837371756520666163696C69736973206D;
        inPKT[900]      = 144'hC384617572697320657520656C656D656E74;
        inPKT[901]      = 144'hC385756D207661726975732E204F72636920;
        inPKT[902]      = 144'hC386766172697573206E61746F7175652070;
        inPKT[903]      = 144'hC387656E617469627573206574206D61676E;
        inPKT[904]      = 144'hC3886973206469732070617274757269656E;
        inPKT[905]      = 144'hC38974206D6F6E7465732C206E6173636574;
        inPKT[906]      = 144'hC38A7572207269646963756C7573206D7573;
        inPKT[907]      = 144'hC38B2E20446F6E6563206469676E69737369;
        inPKT[908]      = 144'hC38C6D206120697073756D20756C74726963;
        inPKT[909]      = 144'hC38D6965732076656E656E617469732E2056;
        inPKT[910]      = 144'hC38E6976616D7573206E756E632076656C69;
        inPKT[911]      = 144'hC38F742C207665686963756C612076697461;
        inPKT[912]      = 144'hC39065206D617373612075742C20636F6E76;
        inPKT[913]      = 144'hC391616C6C697320636F6E73656374657475;
        inPKT[914]      = 144'hC3927220746F72746F722E20517569737175;
        inPKT[915]      = 144'hC3936520616C697175616D2C206E69736C20;
        inPKT[916]      = 144'hC394636F6E67756520626C616E6469742075;
        inPKT[917]      = 144'hC3956C747269636965732C2075726E612074;
        inPKT[918]      = 144'hC3967572706973206D6174746973206D6167;
        inPKT[919]      = 144'hC3976E612C206E6F6E206665726D656E7475;
        inPKT[920]      = 144'hC3986D206475692076656C69742065752071;
        inPKT[921]      = 144'hC39975616D2E0D0A0D0A496E207068617265;
        inPKT[922]      = 144'hC39A7472612076656C697420646F6C6F722C;
        inPKT[923]      = 144'hC39B20766974616520637572737573206F72;
        inPKT[924]      = 144'hC39C63692066696E696275732074696E6369;
        inPKT[925]      = 144'hC39D64756E742E20566976616D7573206964;
        inPKT[926]      = 144'hC39E20746F72746F722072686F6E6375732C;
        inPKT[927]      = 144'hC39F207361676974746973206469616D2065;
        inPKT[928]      = 144'hC3A06765742C207072657469756D206D6175;
        inPKT[929]      = 144'hC3A17269732E2050686173656C6C75732065;
        inPKT[930]      = 144'hC3A26C656D656E74756D20656E696D206665;
        inPKT[931]      = 144'hC3A36C69732E204D6175726973206575206E;
        inPKT[932]      = 144'hC3A465717565206567657420707572757320;
        inPKT[933]      = 144'hC3A568656E64726572697420677261766964;
        inPKT[934]      = 144'hC3A6612E20416C697175616D206C69626572;
        inPKT[935]      = 144'hC3A76F206E6962682C20636F6E76616C6C69;
        inPKT[936]      = 144'hC3A8732061206E69736C2065742C2068656E;
        inPKT[937]      = 144'hC3A964726572697420766573746962756C75;
        inPKT[938]      = 144'hC3AA6D2066656C69732E20446F6E65632065;
        inPKT[939]      = 144'hC3AB7569736D6F64206665726D656E74756D;
        inPKT[940]      = 144'hC3AC2074757270697320657520617563746F;
        inPKT[941]      = 144'hC3AD722E2041656E65616E20626962656E64;
        inPKT[942]      = 144'hC3AE756D2074757270697320696E206F6469;
        inPKT[943]      = 144'hC3AF6F20636F6E76616C6C69732C20766974;
        inPKT[944]      = 144'hC3B0616520766172697573206578206C616F;
        inPKT[945]      = 144'hC3B1726565742E2046757363652076656C20;
        inPKT[946]      = 144'hC3B26D6920766974616520646F6C6F722066;
        inPKT[947]      = 144'hC3B36575676961742076756C707574617465;
        inPKT[948]      = 144'hC3B4206E6563207574206E756E632E204372;
        inPKT[949]      = 144'hC3B5617320646170696275732C20616E7465;
        inPKT[950]      = 144'hC3B6206964207665686963756C6120616C69;
        inPKT[951]      = 144'hC3B77175616D2C20656C69742065726F7320;
        inPKT[952]      = 144'hC3B87361676974746973206D692C206E6F6E;
        inPKT[953]      = 144'hC3B920656C656966656E64206578206E756C;
        inPKT[954]      = 144'hC3BA6C6120656765742076656C69742E2053;
        inPKT[955]      = 144'hC3BB757370656E6469737365206964206469;
        inPKT[956]      = 144'hC3BC616D206475692E2053757370656E6469;
        inPKT[957]      = 144'hC3BD737365207072657469756D206A757374;
        inPKT[958]      = 144'hC3BE6F20736564206E69626820706F727474;
        inPKT[959]      = 144'hC3BF69746F722C2076656C20696E74657264;
        inPKT[960]      = 144'hC3C0756D206D6175726973206D6178696D75;
        inPKT[961]      = 144'hC3C1732E20557420616C697175616D206C61;
        inPKT[962]      = 144'hC3C26375732070757275732C207369742061;
        inPKT[963]      = 144'hC3C36D657420696D70657264696574206E69;
        inPKT[964]      = 144'hC3C4626820666575676961742069642E2049;
        inPKT[965]      = 144'hC3C56E7465676572206C6F72656D206D6175;
        inPKT[966]      = 144'hC3C67269732C207072657469756D206E6F6E;
        inPKT[967]      = 144'hC3C7206E6973692065742C20646170696275;
        inPKT[968]      = 144'hC3C8732066696E69627573206F7263692E0D;
        inPKT[969]      = 144'hC3C90A0D0A566573746962756C756D206961;
        inPKT[970]      = 144'hC3CA63756C69732C206D61676E6120617420;
        inPKT[971]      = 144'hC3CB6D6174746973206D6178696D75732C20;
        inPKT[972]      = 144'hC3CC61726375206572617420646170696275;
        inPKT[973]      = 144'hC3CD73206E756E632C206120766172697573;
        inPKT[974]      = 144'hC3CE206D657475732066656C697320736564;
        inPKT[975]      = 144'hC3CF206F7263692E204E756C6C616D206D69;
        inPKT[976]      = 144'hC3D0206E6962682C20656C656966656E6420;
        inPKT[977]      = 144'hC3D16E656320756C747269636573206E6563;
        inPKT[978]      = 144'hC3D22C20636F6E7365637465747572206163;
        inPKT[979]      = 144'hC3D320656E696D2E20536564206C75637475;
        inPKT[980]      = 144'hC3D4732073656D20717569732074656D706F;
        inPKT[981]      = 144'hC3D57220636F6E6775652E2053757370656E;
        inPKT[982]      = 144'hC3D6646973736520706F74656E74692E2045;
        inPKT[983]      = 144'hC3D77469616D2065676574206C696265726F;
        inPKT[984]      = 144'hC3D82076656C69742E204475697320766573;
        inPKT[985]      = 144'hC3D9746962756C756D20636F6E7365717561;
        inPKT[986]      = 144'hC3DA7420706F7274612E204D617572697320;
        inPKT[987]      = 144'hC3DB706F72747469746F7220747572706973;
        inPKT[988]      = 144'hC3DC20696E206D6173736120616C69717561;
        inPKT[989]      = 144'hC3DD6D20636F6E6775652E204E756C6C6120;
        inPKT[990]      = 144'hC3DE636F6E73656374657475722075726E61;
        inPKT[991]      = 144'hC3DF206D657475732C20696420696163756C;
        inPKT[992]      = 144'hC3E06973206E756E6320756C747269636965;
        inPKT[993]      = 144'hC3E17320656765742E204375726162697475;
        inPKT[994]      = 144'hC3E272206D6175726973206E657175652C20;
        inPKT[995]      = 144'hC3E3626962656E64756D207365642065726F;
        inPKT[996]      = 144'hC3E4732061742C206D6178696D757320756C;
        inPKT[997]      = 144'hC3E5747269636573207475727069732E0D0A;
        inPKT[998]      = 144'hC3E6496E74657264756D206574206D616C65;
        inPKT[999]      = 144'hC3E773756164612066616D65732061632061;
        inPKT[1000]     = 144'hC3E86E746520697073756D207072696D6973;
        inPKT[1001]     = 144'hC3E920696E2066617563696275732E205065;
        inPKT[1002]     = 144'hC3EA6C6C656E74657371756520736F6C6C69;
        inPKT[1003]     = 144'hC3EB6369747564696E20626C616E64697420;
        inPKT[1004]     = 144'hC3EC6665726D656E74756D2E2050656C6C65;
        inPKT[1005]     = 144'hC3ED6E746573717565206E6F6E206C696775;
        inPKT[1006]     = 144'hC3EE6C6120657520657261742076656E656E;
        inPKT[1007]     = 144'hC3EF6174697320657569736D6F642E205065;
        inPKT[1008]     = 144'hC3F06C6C656E74657371756520736F64616C;
        inPKT[1009]     = 144'hC3F1657320766573746962756C756D20636F;
        inPKT[1010]     = 144'hC3F26E76616C6C69732E2050726F696E206D;
        inPKT[1011]     = 144'hC3F36F6C6573746965207072657469756D20;
        inPKT[1012]     = 144'hC3F465726F732076656C2065676573746173;
        inPKT[1013]     = 144'hC3F52E204D6F72626920736F6C6C69636974;
        inPKT[1014]     = 144'hC3F67564696E207075727573206163206665;
        inPKT[1015]     = 144'hC3F7726D656E74756D206D61747469732E20;
        inPKT[1016]     = 144'hC3F84E756E632076656C2074696E63696475;
        inPKT[1017]     = 144'hC3F96E74206C696265726F2E204E756C6C61;
        inPKT[1018]     = 144'hC3FA20616C697175657420697073756D206E;
        inPKT[1019]     = 144'hC3FB6563207175616D20696D706572646965;
        inPKT[1020]     = 144'hC3FC7420696E74657264756D2E2050726165;
        inPKT[1021]     = 144'hC3FD73656E74206C6967756C612066656C69;
        inPKT[1022]     = 144'hC3FE732C20696163756C697320617420616C;
        inPKT[1023]     = 144'hC3FF69717565742061742C20736167697474;
        inPKT[1024]     = 144'hC3006973207175697320656C69742E0D0A51;
        inPKT[1025]     = 144'hC3017569737175652076656C20696D706572;
        inPKT[1026]     = 144'hC30264696574206E6962682E205068617365;
        inPKT[1027]     = 144'hC3036C6C75732072757472756D206469676E;
        inPKT[1028]     = 144'hC304697373696D207269737573206E6F6E20;
        inPKT[1029]     = 144'hC30574696E636964756E742E205665737469;
        inPKT[1030]     = 144'hC30662756C756D206E756E6320697073756D;
        inPKT[1031]     = 144'hC3072C2076656E656E617469732065676574;
        inPKT[1032]     = 144'hC30820706F72746120696E2C20636F6E7365;
        inPKT[1033]     = 144'hC30963746574757220657520657261742E20;
        inPKT[1034]     = 144'hC30A446F6E6563207665686963756C612061;
        inPKT[1035]     = 144'hC30B6E74652076656C2072686F6E63757320;
        inPKT[1036]     = 144'hC30C66617563696275732E2050656C6C656E;
        inPKT[1037]     = 144'hC30D746573717565206A7573746F20746F72;
        inPKT[1038]     = 144'hC30E746F722C20766F6C757470617420696E;
        inPKT[1039]     = 144'hC30F206D61757269732061742C2076617269;
        inPKT[1040]     = 144'hC31075732070686172657472612072697375;
        inPKT[1041]     = 144'hC311732E2051756973717565207574206469;
        inPKT[1042]     = 144'hC312616D2073757363697069742C20736F6C;
        inPKT[1043]     = 144'hC3136C696369747564696E2073617069656E;
        inPKT[1044]     = 144'hC3142065742C20696E74657264756D206C61;
        inPKT[1045]     = 144'hC3156375732E204D6F726269207269737573;
        inPKT[1046]     = 144'hC3162073656D2C2070656C6C656E74657371;
        inPKT[1047]     = 144'hC31775652065742074757270697320696E2C;
        inPKT[1048]     = 144'hC31820626C616E64697420736F6C6C696369;
        inPKT[1049]     = 144'hC319747564696E2073656D2E205365642065;
        inPKT[1050]     = 144'hC31A6666696369747572206C696265726F20;
        inPKT[1051]     = 144'hC31B71756973207072657469756D20707265;
        inPKT[1052]     = 144'hC31C7469756D2E204E756C6C616D20617563;
        inPKT[1053]     = 144'hC31D746F72207361676974746973206C6F72;
        inPKT[1054]     = 144'hC31E656D2C20616320756C74726963657320;
        inPKT[1055]     = 144'hC31F61726375206D6178696D757320656765;
        inPKT[1056]     = 144'hC320742E0D0A566573746962756C756D2076;
        inPKT[1057]     = 144'hC3216F6C7574706174206C6967756C612061;
        inPKT[1058]     = 144'hC3227563746F722073656D20766976657272;
        inPKT[1059]     = 144'hC323612C20756C6C616D636F727065722065;
        inPKT[1060]     = 144'hC3247569736D6F64206E6571756520706F72;
        inPKT[1061]     = 144'hC325747469746F722E2053757370656E6469;
        inPKT[1062]     = 144'hC3267373652076697665727261207363656C;
        inPKT[1063]     = 144'hC32765726973717565206F64696F2072686F;
        inPKT[1064]     = 144'hC3286E63757320766F6C75747061742E2041;
        inPKT[1065]     = 144'hC3296C697175616D206572617420766F6C75;
        inPKT[1066]     = 144'hC32A747061742E2053757370656E64697373;
        inPKT[1067]     = 144'hC32B6520706F74656E74692E20496E206861;
        inPKT[1068]     = 144'hC32C632068616269746173736520706C6174;
        inPKT[1069]     = 144'hC32D65612064696374756D73742E2050726F;
        inPKT[1070]     = 144'hC32E696E207574206E756C6C612075742064;
        inPKT[1071]     = 144'hC32F7569207363656C657269737175652064;
        inPKT[1072]     = 144'hC330696374756D2E20517569737175652073;
        inPKT[1073]     = 144'hC33175736369706974206E69626820706F73;
        inPKT[1074]     = 144'hC33275657265207175616D2076756C707574;
        inPKT[1075]     = 144'hC3336174652C206575206C6163696E696120;
        inPKT[1076]     = 144'hC334616E746520677261766964612E204375;
        inPKT[1077]     = 144'hC33572616269747572206D61737361206C6F;
        inPKT[1078]     = 144'hC33672656D2C206F726E617265206575206D;
        inPKT[1079]     = 144'hC3376F6C6C69732061742C20706861726574;
        inPKT[1080]     = 144'hC3387261206E6563206D617373612E204E75;
        inPKT[1081]     = 144'hC3396C6C612066696E6962757320656C6569;
        inPKT[1082]     = 144'hC33A66656E64206F7263692073697420616D;
        inPKT[1083]     = 144'hC33B657420636F6E73656374657475722E20;
        inPKT[1084]     = 144'hC33C5365642074656D707573207669746165;
        inPKT[1085]     = 144'hC33D2061726375206E6563206665726D656E;
        inPKT[1086]     = 144'hC33E74756D2E2041656E65616E2070656C6C;
        inPKT[1087]     = 144'hC33F656E7465737175652076697461652064;
        inPKT[1088]     = 144'hC3406F6C6F7220696E20616363756D73616E;
        inPKT[1089]     = 144'hC3412E2043726173206469676E697373696D;
        inPKT[1090]     = 144'hC3422076756C707574617465206D6F6C6C69;
        inPKT[1091]     = 144'hC343732E204D617572697320706F72746120;
        inPKT[1092]     = 144'hC34476656E656E617469732072697375732C;
        inPKT[1093]     = 144'hC3452065752074726973746971756520646F;
        inPKT[1094]     = 144'hC3466C6F722072757472756D20696E2E2046;
        inPKT[1095]     = 144'hC3477573636520636F6E64696D656E74756D;
        inPKT[1096]     = 144'hC348206F7263692066656C69732C20736974;
        inPKT[1097]     = 144'hC34920616D657420636F6E76616C6C697320;
        inPKT[1098]     = 144'hC34A6C696265726F2074696E636964756E74;
        inPKT[1099]     = 144'hC34B2061632E0D0A566573746962756C756D;
        inPKT[1100]     = 144'hC34C20696D7065726469657420656C697420;
        inPKT[1101]     = 144'hC34D74656D706F72207175616D2067726176;
        inPKT[1102]     = 144'hC34E6964612C207574206D616C6573756164;
        inPKT[1103]     = 144'hC34F612074656C6C757320696D7065726469;
        inPKT[1104]     = 144'hC35065742E2050686173656C6C7573206F64;
        inPKT[1105]     = 144'hC351696F2073656D2C206D61747469732073;
        inPKT[1106]     = 144'hC352656420756C7472696365732061742C20;
        inPKT[1107]     = 144'hC353766976657272612076656C206475692E;
        inPKT[1108]     = 144'hC354204E756E632075726E61206D65747573;
        inPKT[1109]     = 144'hC3552C206C7563747573206163206D617869;
        inPKT[1110]     = 144'hC3566D757320696E2C20636F6E7365637465;
        inPKT[1111]     = 144'hC357747572206E6F6E206E6973692E204E75;
        inPKT[1112]     = 144'hC3586C6C612073697420616D657420626962;
        inPKT[1113]     = 144'hC359656E64756D2076656C69742E20446F6E;
        inPKT[1114]     = 144'hC35A6563207175697320656E696D206E6F6E;
        inPKT[1115]     = 144'hC35B20726973757320626C616E6469742066;
        inPKT[1116]     = 144'hC35C6163696C697369732071756973206E65;
        inPKT[1117]     = 144'hC35D632072697375732E2043757261626974;
        inPKT[1118]     = 144'hC35E75722065752065737420766974616520;
        inPKT[1119]     = 144'hC35F6C656374757320626C616E6469742061;
        inPKT[1120]     = 144'hC3606C69717565742E20566573746962756C;
        inPKT[1121]     = 144'hC361756D20616E746520697073756D207072;
        inPKT[1122]     = 144'hC362696D697320696E206661756369627573;
        inPKT[1123]     = 144'hC363206F726369206C756374757320657420;
        inPKT[1124]     = 144'hC364756C74726963657320706F7375657265;
        inPKT[1125]     = 144'hC36520637562696C69612043757261653B20;
        inPKT[1126]     = 144'hC366566573746962756C756D206163206469;
        inPKT[1127]     = 144'hC367676E697373696D206E756E632E205175;
        inPKT[1128]     = 144'hC368697371756520696E2073616769747469;
        inPKT[1129]     = 144'hC369732074656C6C75732C2073697420616D;
        inPKT[1130]     = 144'hC36A6574206665726D656E74756D206E6962;
        inPKT[1131]     = 144'hC36B682E0D0A496E206469676E697373696D;
        inPKT[1132]     = 144'hC36C20726973757320766974616520707572;
        inPKT[1133]     = 144'hC36D757320766573746962756C756D2C2061;
        inPKT[1134]     = 144'hC36E7420656C656D656E74756D206E756C6C;
        inPKT[1135]     = 144'hC36F6120706F73756572652E20536564206D;
        inPKT[1136]     = 144'hC3706174746973206E756E63206E6962682E;
        inPKT[1137]     = 144'hC3712053757370656E64697373652070656C;
        inPKT[1138]     = 144'hC3726C656E74657371756520706C61636572;
        inPKT[1139]     = 144'hC3736174207363656C657269737175652E20;
        inPKT[1140]     = 144'hC37441656E65616E2066657567696174206D;
        inPKT[1141]     = 144'hC375617572697320696420636F6E67756520;
        inPKT[1142]     = 144'hC3766C6163696E69612E20457469616D2073;
        inPKT[1143]     = 144'hC37775736369706974206C6967756C612074;
        inPKT[1144]     = 144'hC378656C6C75732C206120636F6E67756520;
        inPKT[1145]     = 144'hC3796C656374757320616C697175616D2076;
        inPKT[1146]     = 144'hC37A65686963756C612E2053757370656E64;
        inPKT[1147]     = 144'hC37B69737365206567657420616E74652076;
        inPKT[1148]     = 144'hC37C656C20656E696D206D616C6573756164;
        inPKT[1149]     = 144'hC37D6120766976657272612E2050726F696E;
        inPKT[1150]     = 144'hC37E2074696E636964756E74206172637520;
        inPKT[1151]     = 144'hC37F656765742076756C7075746174652061;
        inPKT[1152]     = 144'hC3806363756D73616E2E20496E2076697461;
        inPKT[1153]     = 144'hC38165206469616D206E6962682E204D6F72;
        inPKT[1154]     = 144'hC3826269206D6178696D75732066656C6973;
        inPKT[1155]     = 144'hC38320696420636F6E736563746574757220;
        inPKT[1156]     = 144'hC384616C697175616D2E204E756C6C612066;
        inPKT[1157]     = 144'hC3856163696C6973692E0D0A566573746962;
        inPKT[1158]     = 144'hC386756C756D20766573746962756C756D20;
        inPKT[1159]     = 144'hC38765666669636974757220746F72746F72;
        inPKT[1160]     = 144'hC3882073697420616D657420666163696C69;
        inPKT[1161]     = 144'hC3897369732E204D616563656E6173206E6F;
        inPKT[1162]     = 144'hC38A6E2074656C6C7573206F7263692E2050;
        inPKT[1163]     = 144'hC38B686173656C6C7573206E6F6E206C7563;
        inPKT[1164]     = 144'hC38C747573206A7573746F2C206174207375;
        inPKT[1165]     = 144'hC38D7363697069742074656C6C75732E2046;
        inPKT[1166]     = 144'hC38E757363652068656E647265726974206E;
        inPKT[1167]     = 144'hC38F6563206E6962682076656C2063757273;
        inPKT[1168]     = 144'hC39075732E2053757370656E646973736520;
        inPKT[1169]     = 144'hC391706F74656E74692E2044756973206C69;
        inPKT[1170]     = 144'hC39267756C612066656C69732C2065666669;
        inPKT[1171]     = 144'hC39363697475722065742076656C69742061;
        inPKT[1172]     = 144'hC394742C20666163696C6973697320636F6E;
        inPKT[1173]     = 144'hC39576616C6C6973206A7573746F2E204E75;
        inPKT[1174]     = 144'hC3966C6C616D206C6F626F72746973207065;
        inPKT[1175]     = 144'hC3976C6C656E74657371756520736F6C6C69;
        inPKT[1176]     = 144'hC3986369747564696E2E204E616D20736974;
        inPKT[1177]     = 144'hC39920616D657420646F6C6F722073697420;
        inPKT[1178]     = 144'hC39A616D6574206C656374757320696D7065;
        inPKT[1179]     = 144'hC39B726469657420636F6E7365717561742E;
        inPKT[1180]     = 144'hC39C20416C697175616D206C756374757320;
        inPKT[1181]     = 144'hC39D7363656C657269737175652070757275;
        inPKT[1182]     = 144'hC39E732C206964206672696E67696C6C6120;
        inPKT[1183]     = 144'hC39F73656D20766F6C75747061742061632E;
        inPKT[1184]     = 144'hC3A0205365642074656D706F722C20656E69;
        inPKT[1185]     = 144'hC3A16D206567657420657569736D6F642066;
        inPKT[1186]     = 144'hC3A26163696C697369732C206E6973692065;
        inPKT[1187]     = 144'hC3A3782073656D70657220697073756D2C20;
        inPKT[1188]     = 144'hC3A4696E207361676974746973206F726369;
        inPKT[1189]     = 144'hC3A5207175616D20696E206C65637475732E;
        inPKT[1190]     = 144'hC3A620557420766974616520656C6974206C;
        inPKT[1191]     = 144'hC3A76967756C612E204E756E632065676573;
        inPKT[1192]     = 144'hC3A87461732C206D69207669746165206961;
        inPKT[1193]     = 144'hC3A963756C6973206D61747469732C206475;
        inPKT[1194]     = 144'hC3AA69206E69626820656C656966656E6420;
        inPKT[1195]     = 144'hC3AB6E69736C2C206567657420706F727461;
        inPKT[1196]     = 144'hC3AC206C696265726F206175677565207175;
        inPKT[1197]     = 144'hC3AD697320656E696D2E2053656420736974;
        inPKT[1198]     = 144'hC3AE20616D65742070756C76696E61722065;
        inPKT[1199]     = 144'hC3AF782C2076656C2070656C6C656E746573;
        inPKT[1200]     = 144'hC3B0717565206C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
