`include "SIMON_defintions.svh"

module test_SIMON_64128_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 1201
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 144'hE4001B1A1918131211100B0A090803020100;
        inPKT[1]        = 144'hC401656B696C20646E75656B696C20646E75;
        inPKT[2]        = 144'hC4024C6F72656D20697073756D20646F6C6F;
        inPKT[3]        = 144'hC403722073697420616D65742C20636F6E73;
        inPKT[4]        = 144'hC40465637465747572206164697069736369;
        inPKT[5]        = 144'hC4056E6720656C69742E2043757261626974;
        inPKT[6]        = 144'hC406757220756C6C616D636F727065722074;
        inPKT[7]        = 144'hC407656D707573206E6973692C2065742070;
        inPKT[8]        = 144'hC4086F73756572652075726E612E2041656E;
        inPKT[9]        = 144'hC40965616E20736564206772617669646120;
        inPKT[10]       = 144'hC40A6C616375732E204E756C6C6120666163;
        inPKT[11]       = 144'hC40B696C6973692E204E756C6C612074656D;
        inPKT[12]       = 144'hC40C707573206F726369207175697320656C;
        inPKT[13]       = 144'hC40D697420666575676961742C2076656C20;
        inPKT[14]       = 144'hC40E73656D706572206C656F20696D706572;
        inPKT[15]       = 144'hC40F646965742E204D616563656E61732065;
        inPKT[16]       = 144'hC41074206E756E6320696E206E6962682066;
        inPKT[17]       = 144'hC4116163696C6973697320636F6E76616C6C;
        inPKT[18]       = 144'hC41269732E2053656420636F6E6775652068;
        inPKT[19]       = 144'hC413656E64726572697420696163756C6973;
        inPKT[20]       = 144'hC4142E20566976616D757320766568696375;
        inPKT[21]       = 144'hC4156C61206C7563747573206573742C2076;
        inPKT[22]       = 144'hC41669746165207375736369706974206E69;
        inPKT[23]       = 144'hC417736C20706F72747469746F722061632E;
        inPKT[24]       = 144'hC4180D0A0D0A446F6E6563206D6F6C657374;
        inPKT[25]       = 144'hC41969652073617069656E2069642076756C;
        inPKT[26]       = 144'hC41A70757461746520766573746962756C75;
        inPKT[27]       = 144'hC41B6D2E204E756C6C6120696E206C696775;
        inPKT[28]       = 144'hC41C6C61206672696E67696C6C612C20756C;
        inPKT[29]       = 144'hC41D6C616D636F727065722075726E612065;
        inPKT[30]       = 144'hC41E742C20706F72747469746F72206C6563;
        inPKT[31]       = 144'hC41F7475732E205175697371756520626C61;
        inPKT[32]       = 144'hC4206E646974206575206D61757269732061;
        inPKT[33]       = 144'hC421632068656E6472657269742E204E756C;
        inPKT[34]       = 144'hC4226C612076656E656E617469732C206D65;
        inPKT[35]       = 144'hC423747573206574206C7563747573206672;
        inPKT[36]       = 144'hC424696E67696C6C612C206E696268207665;
        inPKT[37]       = 144'hC4256C697420756C6C616D636F7270657220;
        inPKT[38]       = 144'hC4266469616D2C2065676574206566666963;
        inPKT[39]       = 144'hC4276974757220697073756D207475727069;
        inPKT[40]       = 144'hC42873206174206E6962682E205574206567;
        inPKT[41]       = 144'hC4296574207072657469756D2065726F732C;
        inPKT[42]       = 144'hC42A20656765742064696374756D206C6163;
        inPKT[43]       = 144'hC42B75732E204D616563656E617320757420;
        inPKT[44]       = 144'hC42C656E696D2065782E2041656E65616E20;
        inPKT[45]       = 144'hC42D76697461652073656D7065722066656C;
        inPKT[46]       = 144'hC42E69732C2073656420756C747269636965;
        inPKT[47]       = 144'hC42F732072697375732E20446F6E65632063;
        inPKT[48]       = 144'hC4306F6E7365637465747572206D69206E69;
        inPKT[49]       = 144'hC431736C2C20617420637572737573206970;
        inPKT[50]       = 144'hC43273756D206772617669646120612E2050;
        inPKT[51]       = 144'hC433686173656C6C75732073697420616D65;
        inPKT[52]       = 144'hC43474206D61676E612076656C2069707375;
        inPKT[53]       = 144'hC4356D206567657374617320706F7274612E;
        inPKT[54]       = 144'hC43620566976616D7573206C756374757320;
        inPKT[55]       = 144'hC437656E696D20656765742074656D706F72;
        inPKT[56]       = 144'hC4382073616769747469732E20416C697175;
        inPKT[57]       = 144'hC439616D20626962656E64756D2073656D20;
        inPKT[58]       = 144'hC43A6120636F6E7365637465747572206566;
        inPKT[59]       = 144'hC43B666963697475722E20446F6E65632073;
        inPKT[60]       = 144'hC43C63656C6572697371756520616C697175;
        inPKT[61]       = 144'hC43D616D206375727375732E204375726162;
        inPKT[62]       = 144'hC43E697475722073697420616D6574206269;
        inPKT[63]       = 144'hC43F62656E64756D20656C69742E20536564;
        inPKT[64]       = 144'hC440206469616D206A7573746F2C20696163;
        inPKT[65]       = 144'hC441756C69732071756973206E756C6C6120;
        inPKT[66]       = 144'hC44276697461652C20616C697175616D2065;
        inPKT[67]       = 144'hC4437569736D6F642066656C69732E0D0A0D;
        inPKT[68]       = 144'hC4440A50726F696E20646170696275732C20;
        inPKT[69]       = 144'hC4456469616D2076756C7075746174652066;
        inPKT[70]       = 144'hC44672696E67696C6C61206D616C65737561;
        inPKT[71]       = 144'hC44764612C206A7573746F20707572757320;
        inPKT[72]       = 144'hC448636F6D6D6F646F20646F6C6F722C2075;
        inPKT[73]       = 144'hC449742064696374756D2065726174206E75;
        inPKT[74]       = 144'hC44A6E632072757472756D2075726E612E20;
        inPKT[75]       = 144'hC44B4E756C6C612067726176696461207572;
        inPKT[76]       = 144'hC44C6E6120766974616520696D7065726469;
        inPKT[77]       = 144'hC44D6574206C616F726565742E2050656C6C;
        inPKT[78]       = 144'hC44E656E7465737175652072686F6E637573;
        inPKT[79]       = 144'hC44F20626962656E64756D206E6962682C20;
        inPKT[80]       = 144'hC4506964206D6F6C6C6973206469616D2073;
        inPKT[81]       = 144'hC451757363697069742061632E2050656C6C;
        inPKT[82]       = 144'hC452656E7465737175652076656C20696163;
        inPKT[83]       = 144'hC453756C6973206475692E204D6F72626920;
        inPKT[84]       = 144'hC454617420616C6971756574206D61737361;
        inPKT[85]       = 144'hC4552E2050726F696E207669746165206F72;
        inPKT[86]       = 144'hC4566E617265206F64696F2C206575207675;
        inPKT[87]       = 144'hC4576C70757461746520697073756D2E2050;
        inPKT[88]       = 144'hC458726F696E206C6F626F727469732C2073;
        inPKT[89]       = 144'hC459656D206E656320657569736D6F642074;
        inPKT[90]       = 144'hC45A696E636964756E742C20617567756520;
        inPKT[91]       = 144'hC45B6D6175726973207363656C6572697371;
        inPKT[92]       = 144'hC45C7565206D61676E612C20657420706F73;
        inPKT[93]       = 144'hC45D75657265206D69206E69736C206E6563;
        inPKT[94]       = 144'hC45E206E6973692E20467573636520656C69;
        inPKT[95]       = 144'hC45F74206E657175652C2076617269757320;
        inPKT[96]       = 144'hC4606574206672696E67696C6C6120766974;
        inPKT[97]       = 144'hC46161652C207661726975732076656C206E;
        inPKT[98]       = 144'hC462657175652E204E756C6C612065742074;
        inPKT[99]       = 144'hC463656D707573206A7573746F2E204D6F72;
        inPKT[100]      = 144'hC464626920756C6C616D636F727065722073;
        inPKT[101]      = 144'hC4657573636970697420636F6E6775652E20;
        inPKT[102]      = 144'hC46653656420656C656966656E64206F6469;
        inPKT[103]      = 144'hC4676F206163207375736369706974206469;
        inPKT[104]      = 144'hC468676E697373696D2E2051756973717565;
        inPKT[105]      = 144'hC46920616E746520656E696D2C20626C616E;
        inPKT[106]      = 144'hC46A64697420696E20636F6E736571756174;
        inPKT[107]      = 144'hC46B2061632C20696E74657264756D207669;
        inPKT[108]      = 144'hC46C7461652070757275732E204D61757269;
        inPKT[109]      = 144'hC46D7320657569736D6F6420706F73756572;
        inPKT[110]      = 144'hC46E65206C65637475732E20566976616D75;
        inPKT[111]      = 144'hC46F7320696E74657264756D207175616D20;
        inPKT[112]      = 144'hC47065752073656D70657220666175636962;
        inPKT[113]      = 144'hC47175732E0D0A0D0A496E206D6F6C657374;
        inPKT[114]      = 144'hC4726965206E756C6C6120616E74652C2061;
        inPKT[115]      = 144'hC4736320696E74657264756D206D61676E61;
        inPKT[116]      = 144'hC47420636F6E64696D656E74756D20636F6E;
        inPKT[117]      = 144'hC47564696D656E74756D2E20447569732075;
        inPKT[118]      = 144'hC4766C7472696369657320736F64616C6573;
        inPKT[119]      = 144'hC477206E756C6C612C2073697420616D6574;
        inPKT[120]      = 144'hC47820756C6C616D636F72706572206F6469;
        inPKT[121]      = 144'hC4796F207072657469756D206E65632E2046;
        inPKT[122]      = 144'hC47A75736365207365642072697375732070;
        inPKT[123]      = 144'hC47B656C6C656E7465737175652C20636F6E;
        inPKT[124]      = 144'hC47C76616C6C69732073656D20656765742C;
        inPKT[125]      = 144'hC47D2068656E64726572697420657261742E;
        inPKT[126]      = 144'hC47E204D6F72626920736F64616C65732076;
        inPKT[127]      = 144'hC47F65686963756C61206C6F626F72746973;
        inPKT[128]      = 144'hC4802E2041656E65616E206120746F72746F;
        inPKT[129]      = 144'hC48172206375727375732C207363656C6572;
        inPKT[130]      = 144'hC4826973717565206C6967756C6120706F72;
        inPKT[131]      = 144'hC483747469746F722C206567657374617320;
        inPKT[132]      = 144'hC48465726F732E20447569732074696E6369;
        inPKT[133]      = 144'hC48564756E7420746F72746F722069642070;
        inPKT[134]      = 144'hC4866F737565726520677261766964612E20;
        inPKT[135]      = 144'hC487496E20636F6E76616C6C6973206D6920;
        inPKT[136]      = 144'hC488696420697073756D206D616C65737561;
        inPKT[137]      = 144'hC48964612C2075742064696374756D206572;
        inPKT[138]      = 144'hC48A6F7320696D706572646965742E205072;
        inPKT[139]      = 144'hC48B6F696E20756C6C616D636F727065722C;
        inPKT[140]      = 144'hC48C206D6175726973206964207661726975;
        inPKT[141]      = 144'hC48D7320636F6E6775652C2065726F732073;
        inPKT[142]      = 144'hC48E617069656E2072686F6E637573206D69;
        inPKT[143]      = 144'hC48F2C20617420617563746F72206E657175;
        inPKT[144]      = 144'hC490652061726375206C616F726565742064;
        inPKT[145]      = 144'hC49169616D2E0D0A0D0A467573636520706F;
        inPKT[146]      = 144'hC49272747469746F72206C696265726F2061;
        inPKT[147]      = 144'hC4937263752C206C6163696E69612068656E;
        inPKT[148]      = 144'hC494647265726974206469616D20636F6E76;
        inPKT[149]      = 144'hC495616C6C6973207365642E205068617365;
        inPKT[150]      = 144'hC4966C6C7573206E6F6E2074757270697320;
        inPKT[151]      = 144'hC49770686172657472612C20756C6C616D63;
        inPKT[152]      = 144'hC4986F72706572206E657175652076656C2C;
        inPKT[153]      = 144'hC49920736F6C6C696369747564696E207665;
        inPKT[154]      = 144'hC49A6C69742E2050656C6C656E7465737175;
        inPKT[155]      = 144'hC49B65206861626974616E74206D6F726269;
        inPKT[156]      = 144'hC49C207472697374697175652073656E6563;
        inPKT[157]      = 144'hC49D747573206574206E6574757320657420;
        inPKT[158]      = 144'hC49E6D616C6573756164612066616D657320;
        inPKT[159]      = 144'hC49F61632074757270697320656765737461;
        inPKT[160]      = 144'hC4A0732E204E616D206E6563207361706965;
        inPKT[161]      = 144'hC4A16E206D6F6C65737469652C2064696374;
        inPKT[162]      = 144'hC4A2756D206D6173736120656765742C2065;
        inPKT[163]      = 144'hC4A3676573746173206F64696F2E20457469;
        inPKT[164]      = 144'hC4A4616D20617263752073617069656E2C20;
        inPKT[165]      = 144'hC4A57072657469756D2061206D6F6C6C6973;
        inPKT[166]      = 144'hC4A620612C2076756C707574617465206E6F;
        inPKT[167]      = 144'hC4A76E20657261742E205574207669746165;
        inPKT[168]      = 144'hC4A8206E696268206C6F626F72746973206C;
        inPKT[169]      = 144'hC4A965637475732066617563696275732070;
        inPKT[170]      = 144'hC4AA6F7274612065752073697420616D6574;
        inPKT[171]      = 144'hC4AB206E69736C2E204D6F72626920706F72;
        inPKT[172]      = 144'hC4AC747469746F722076656C697420657520;
        inPKT[173]      = 144'hC4AD646F6C6F72206C616F726565742C2073;
        inPKT[174]      = 144'hC4AE697420616D657420696D706572646965;
        inPKT[175]      = 144'hC4AF7420656E696D20736F64616C65732E20;
        inPKT[176]      = 144'hC4B04E756C6C616D20756C6C616D636F7270;
        inPKT[177]      = 144'hC4B16572207475727069732061742070656C;
        inPKT[178]      = 144'hC4B26C656E74657371756520766172697573;
        inPKT[179]      = 144'hC4B32E20566976616D757320657520696D70;
        inPKT[180]      = 144'hC4B4657264696574206E657175652E205365;
        inPKT[181]      = 144'hC4B564207175697320617563746F7220616E;
        inPKT[182]      = 144'hC4B674652E204D61757269732073656D7065;
        inPKT[183]      = 144'hC4B77220697073756D207365642064756920;
        inPKT[184]      = 144'hC4B8706F73756572652C20617420616C6971;
        inPKT[185]      = 144'hC4B975616D206D6574757320656C65696665;
        inPKT[186]      = 144'hC4BA6E642E204E756C6C616D207472697374;
        inPKT[187]      = 144'hC4BB6971756520656C656966656E64206572;
        inPKT[188]      = 144'hC4BC6F732C2065676574206665726D656E74;
        inPKT[189]      = 144'hC4BD756D20697073756D20656C656D656E74;
        inPKT[190]      = 144'hC4BE756D206E65632E0D0A0D0A50656C6C65;
        inPKT[191]      = 144'hC4BF6E7465737175652068656E6472657269;
        inPKT[192]      = 144'hC4C07420626962656E64756D206C6967756C;
        inPKT[193]      = 144'hC4C1612C20657420736F64616C6573206D61;
        inPKT[194]      = 144'hC4C2676E61206461706962757320696E2E20;
        inPKT[195]      = 144'hC4C3496E20616C697175657420746F72746F;
        inPKT[196]      = 144'hC4C472206567657420636F6E736563746574;
        inPKT[197]      = 144'hC4C5757220636F6E73656374657475722E20;
        inPKT[198]      = 144'hC4C651756973717565207472697374697175;
        inPKT[199]      = 144'hC4C76520726973757320657261742C206574;
        inPKT[200]      = 144'hC4C820616C697175657420656C697420616C;
        inPKT[201]      = 144'hC4C969717565742065752E20496E74656765;
        inPKT[202]      = 144'hC4CA72206E6F6E206D61676E6120696E2066;
        inPKT[203]      = 144'hC4CB656C697320706F72747469746F722073;
        inPKT[204]      = 144'hC4CC616769747469732E2051756973717565;
        inPKT[205]      = 144'hC4CD2076697665727261206F726369206163;
        inPKT[206]      = 144'hC4CE2072757472756D206C616F726565742E;
        inPKT[207]      = 144'hC4CF2041656E65616E20636F6E76616C6C69;
        inPKT[208]      = 144'hC4D0732064696374756D207475727069732C;
        inPKT[209]      = 144'hC4D12065742066696E696275732073617069;
        inPKT[210]      = 144'hC4D2656E20636F6E67756520696E2E205365;
        inPKT[211]      = 144'hC4D36420612065726174206F726E6172652C;
        inPKT[212]      = 144'hC4D4206D6F6C6C6973206E69736C2061632C;
        inPKT[213]      = 144'hC4D5206469676E697373696D206E65717565;
        inPKT[214]      = 144'hC4D62E2051756973717565206D616C657375;
        inPKT[215]      = 144'hC4D761646120706F73756572652074757270;
        inPKT[216]      = 144'hC4D8697320657520756C6C616D636F727065;
        inPKT[217]      = 144'hC4D9722E20446F6E65632076697665727261;
        inPKT[218]      = 144'hC4DA20626962656E64756D206E756E632C20;
        inPKT[219]      = 144'hC4DB64696374756D20696D70657264696574;
        inPKT[220]      = 144'hC4DC206E65717565206D6178696D75732069;
        inPKT[221]      = 144'hC4DD6E2E20446F6E656320757420756C7472;
        inPKT[222]      = 144'hC4DE6963657320646F6C6F722E2056697661;
        inPKT[223]      = 144'hC4DF6D757320736564206175677565207072;
        inPKT[224]      = 144'hC4E0657469756D2C20766F6C757470617420;
        inPKT[225]      = 144'hC4E1657261742061632C20706F7274612064;
        inPKT[226]      = 144'hC4E269616D2E204D617572697320696E2070;
        inPKT[227]      = 144'hC4E37572757320756C747269636965732C20;
        inPKT[228]      = 144'hC4E47375736369706974206469616D207365;
        inPKT[229]      = 144'hC4E5642C2074696E636964756E7420656E69;
        inPKT[230]      = 144'hC4E66D2E20446F6E6563207175697320706F;
        inPKT[231]      = 144'hC4E77375657265206E6962682E20496E2068;
        inPKT[232]      = 144'hC4E861632068616269746173736520706C61;
        inPKT[233]      = 144'hC4E97465612064696374756D73742E0D0A0D;
        inPKT[234]      = 144'hC4EA0A4D6F726269206F726E617265206A75;
        inPKT[235]      = 144'hC4EB73746F206174207175616D2066617563;
        inPKT[236]      = 144'hC4EC696275732C2073697420616D6574206D;
        inPKT[237]      = 144'hC4ED6F6C6573746965206C656F2063757273;
        inPKT[238]      = 144'hC4EE75732E204D6175726973206C616F7265;
        inPKT[239]      = 144'hC4EF657420616E74652061206D6574757320;
        inPKT[240]      = 144'hC4F065666669636974757220766172697573;
        inPKT[241]      = 144'hC4F12E205365642076656C206F7263692073;
        inPKT[242]      = 144'hC4F261676974746973206E756E6320626C61;
        inPKT[243]      = 144'hC4F36E64697420636F6E7365717561742E20;
        inPKT[244]      = 144'hC4F45072616573656E74206D616C65737561;
        inPKT[245]      = 144'hC4F56461206E657175652071756973206469;
        inPKT[246]      = 144'hC4F66374756D206469676E697373696D2E20;
        inPKT[247]      = 144'hC4F7446F6E656320666163696C6973697320;
        inPKT[248]      = 144'hC4F873697420616D65742076656C69742065;
        inPKT[249]      = 144'hC4F975206C6F626F727469732E204E756C6C;
        inPKT[250]      = 144'hC4FA616D20626C616E64697420656C656D65;
        inPKT[251]      = 144'hC4FB6E74756D206D61757269732C20766974;
        inPKT[252]      = 144'hC4FC616520656C656D656E74756D20646F6C;
        inPKT[253]      = 144'hC4FD6F722068656E64726572697420766974;
        inPKT[254]      = 144'hC4FE61652E204675736365206D6F6C657374;
        inPKT[255]      = 144'hC4FF69652C20656C697420757420616C6971;
        inPKT[256]      = 144'hC40075657420766F6C75747061742C206E65;
        inPKT[257]      = 144'hC4017175652076656C697420707265746975;
        inPKT[258]      = 144'hC4026D2061756775652C206672696E67696C;
        inPKT[259]      = 144'hC4036C6120636F6E64696D656E74756D206A;
        inPKT[260]      = 144'hC4047573746F2073617069656E2061206A75;
        inPKT[261]      = 144'hC40573746F2E2050686173656C6C75732071;
        inPKT[262]      = 144'hC40675697320617563746F72206C6F72656D;
        inPKT[263]      = 144'hC4072C20696E20616C697175616D206E756E;
        inPKT[264]      = 144'hC408632E20557420656C656966656E642061;
        inPKT[265]      = 144'hC4096E7465206574206E697369206D6F6C65;
        inPKT[266]      = 144'hC40A7374696520636F6E76616C6C69732069;
        inPKT[267]      = 144'hC40B642065742073656D2E20536564206163;
        inPKT[268]      = 144'hC40C20626962656E64756D20617263752E20;
        inPKT[269]      = 144'hC40D467573636520766573746962756C756D;
        inPKT[270]      = 144'hC40E206E756E6320656765742074656C6C75;
        inPKT[271]      = 144'hC40F73206665726D656E74756D2C206E6563;
        inPKT[272]      = 144'hC4102072686F6E637573206D617373612063;
        inPKT[273]      = 144'hC4116F6D6D6F646F2E204D616563656E6173;
        inPKT[274]      = 144'hC412206964206E756E63206E6F6E20657820;
        inPKT[275]      = 144'hC413766573746962756C756D206F726E6172;
        inPKT[276]      = 144'hC41465207574206E65632065726F732E2041;
        inPKT[277]      = 144'hC4156C697175616D20656666696369747572;
        inPKT[278]      = 144'hC41620636F6D6D6F646F206469616D206964;
        inPKT[279]      = 144'hC417206C6F626F727469732E205365642061;
        inPKT[280]      = 144'hC418632074656D706F72206C65637475732E;
        inPKT[281]      = 144'hC419204E756E6320656C656D656E74756D20;
        inPKT[282]      = 144'hC41A7574206C65637475732061632074696E;
        inPKT[283]      = 144'hC41B636964756E742E20557420696163756C;
        inPKT[284]      = 144'hC41C6973206E756C6C612071756973206578;
        inPKT[285]      = 144'hC41D20656C656D656E74756D2C20616C6971;
        inPKT[286]      = 144'hC41E7565742073656D706572206D61676E61;
        inPKT[287]      = 144'hC41F20656C656966656E642E0D0A0D0A4375;
        inPKT[288]      = 144'hC4207261626974757220746F72746F72206E;
        inPKT[289]      = 144'hC42169736C2C20756C747269636965732069;
        inPKT[290]      = 144'hC4226E206E657175652061632C2061636375;
        inPKT[291]      = 144'hC4236D73616E20636F6E736571756174206D;
        inPKT[292]      = 144'hC424657475732E204D616563656E6173206D;
        inPKT[293]      = 144'hC425617373612073617069656E2C206D6174;
        inPKT[294]      = 144'hC42674697320696E2076656E656E61746973;
        inPKT[295]      = 144'hC4272073697420616D65742C20617563746F;
        inPKT[296]      = 144'hC428722073697420616D657420656E696D2E;
        inPKT[297]      = 144'hC429204E756E63207669746165206D657475;
        inPKT[298]      = 144'hC42A7320636F6D6D6F646F2C206D61747469;
        inPKT[299]      = 144'hC42B73206D617373612073697420616D6574;
        inPKT[300]      = 144'hC42C2C20766172697573206C6F72656D2E20;
        inPKT[301]      = 144'hC42D4E756E6320696E20656C697420656C69;
        inPKT[302]      = 144'hC42E742E204E756E63206F726E6172652063;
        inPKT[303]      = 144'hC42F6F6E7365637465747572206D61676E61;
        inPKT[304]      = 144'hC4302C2073697420616D657420706F727474;
        inPKT[305]      = 144'hC43169746F7220617263752072686F6E6375;
        inPKT[306]      = 144'hC432732065752E2053757370656E64697373;
        inPKT[307]      = 144'hC43365207363656C6572697371756520756C;
        inPKT[308]      = 144'hC43474726963696573206578206120616C69;
        inPKT[309]      = 144'hC4357175616D2E2053757370656E64697373;
        inPKT[310]      = 144'hC436652072757472756D20736F6C6C696369;
        inPKT[311]      = 144'hC437747564696E206E756E632C206E6F6E20;
        inPKT[312]      = 144'hC438636F6E76616C6C697320747572706973;
        inPKT[313]      = 144'hC439206C616F726565742073697420616D65;
        inPKT[314]      = 144'hC43A742E2041656E65616E20612066696E69;
        inPKT[315]      = 144'hC43B627573206D61757269732C2071756973;
        inPKT[316]      = 144'hC43C20637572737573206E756E632E20496E;
        inPKT[317]      = 144'hC43D2066657567696174206475692076656C;
        inPKT[318]      = 144'hC43E2075726E612073656D70657220666175;
        inPKT[319]      = 144'hC43F63696275732E204D617572697320756C;
        inPKT[320]      = 144'hC44074726963696573206174207475727069;
        inPKT[321]      = 144'hC4417320656765742070656C6C656E746573;
        inPKT[322]      = 144'hC4427175652E205072616573656E74207369;
        inPKT[323]      = 144'hC4437420616D6574206C6967756C6120636F;
        inPKT[324]      = 144'hC4446E76616C6C69732C20656C656D656E74;
        inPKT[325]      = 144'hC445756D206E756C6C6120756C6C616D636F;
        inPKT[326]      = 144'hC446727065722C20616C697175616D207572;
        inPKT[327]      = 144'hC4476E612E20457469616D207175616D2065;
        inPKT[328]      = 144'hC4486C69742C20706F737565726520757420;
        inPKT[329]      = 144'hC4497175616D20656765742C2066696E6962;
        inPKT[330]      = 144'hC44A757320736F6C6C696369747564696E20;
        inPKT[331]      = 144'hC44B6E756C6C612E20496E20737573636970;
        inPKT[332]      = 144'hC44C697420656E696D2065742065726F7320;
        inPKT[333]      = 144'hC44D66696E696275732C207574207363656C;
        inPKT[334]      = 144'hC44E657269737175652074656C6C75732066;
        inPKT[335]      = 144'hC44F6575676961742E204375726162697475;
        inPKT[336]      = 144'hC45072206E6F6E206D617373612076617269;
        inPKT[337]      = 144'hC451757320646F6C6F722067726176696461;
        inPKT[338]      = 144'hC45220656C656D656E74756D207175697320;
        inPKT[339]      = 144'hC45375742066656C69732E2050686173656C;
        inPKT[340]      = 144'hC4546C757320657569736D6F642069707375;
        inPKT[341]      = 144'hC4556D20656765742076656C6974206C6F62;
        inPKT[342]      = 144'hC4566F727469732C206567657420706F7274;
        inPKT[343]      = 144'hC45761206D61757269732074656D7075732E;
        inPKT[344]      = 144'hC4582053656420696D706572646965742076;
        inPKT[345]      = 144'hC4596F6C75747061742074656C6C75732065;
        inPKT[346]      = 144'hC45A752074696E636964756E742E0D0A0D0A;
        inPKT[347]      = 144'hC45B55742076656C206D69206174206D6574;
        inPKT[348]      = 144'hC45C7573206672696E67696C6C6120677261;
        inPKT[349]      = 144'hC45D766964612E205072616573656E742065;
        inPKT[350]      = 144'hC45E726F73206E6962682C20637572737573;
        inPKT[351]      = 144'hC45F20656765737461732074696E63696475;
        inPKT[352]      = 144'hC4606E7420736F64616C65732C207363656C;
        inPKT[353]      = 144'hC46165726973717565206E65632066656C69;
        inPKT[354]      = 144'hC462732E20496E746567657220696D706572;
        inPKT[355]      = 144'hC46364696574206D616C657375616461206E;
        inPKT[356]      = 144'hC46469736C20616C69717565742076656E65;
        inPKT[357]      = 144'hC4656E617469732E20496E74656765722073;
        inPKT[358]      = 144'hC466656420706F72747469746F7220697073;
        inPKT[359]      = 144'hC467756D2E20496E746567657220636F6D6D;
        inPKT[360]      = 144'hC4686F646F206665756769617420746F7274;
        inPKT[361]      = 144'hC4696F722C206575206C6F626F7274697320;
        inPKT[362]      = 144'hC46A617567756520656C656D656E74756D20;
        inPKT[363]      = 144'hC46B73697420616D65742E20446F6E656320;
        inPKT[364]      = 144'hC46C766573746962756C756D206C6967756C;
        inPKT[365]      = 144'hC46D612061756775652C2065742066696E69;
        inPKT[366]      = 144'hC46E627573206172637520706F7274612069;
        inPKT[367]      = 144'hC46F6E2E204E756C6C612073656D2074656C;
        inPKT[368]      = 144'hC4706C75732C20756C6C616D636F72706572;
        inPKT[369]      = 144'hC4712061742063757273757320612C20706F;
        inPKT[370]      = 144'hC4727274612073697420616D6574206D6167;
        inPKT[371]      = 144'hC4736E612E204E756E632076697461652069;
        inPKT[372]      = 144'hC4746D706572646965742070757275732C20;
        inPKT[373]      = 144'hC4756E656320736F6C6C696369747564696E;
        inPKT[374]      = 144'hC4762074656C6C75732E20416C697175616D;
        inPKT[375]      = 144'hC477206572617420766F6C75747061742E20;
        inPKT[376]      = 144'hC478536564206964206D61676E6120636F6D;
        inPKT[377]      = 144'hC4796D6F646F2C206C75637475732076656C;
        inPKT[378]      = 144'hC47A697420717569732C20657569736D6F64;
        inPKT[379]      = 144'hC47B20656E696D2E20496E7465676572206D;
        inPKT[380]      = 144'hC47C617474697320736F64616C6573206665;
        inPKT[381]      = 144'hC47D726D656E74756D2E2051756973717565;
        inPKT[382]      = 144'hC47E20736564206672696E67696C6C61206C;
        inPKT[383]      = 144'hC47F6F72656D2E2043726173207665686963;
        inPKT[384]      = 144'hC480756C612074656D707573207361706965;
        inPKT[385]      = 144'hC4816E20757420636F6E6775652E20447569;
        inPKT[386]      = 144'hC482732073617069656E20656E696D2C2070;
        inPKT[387]      = 144'hC4836F727461206E6563206C656F2069642C;
        inPKT[388]      = 144'hC4842065666669636974757220706F737565;
        inPKT[389]      = 144'hC4857265206C696265726F2E204E756C6C61;
        inPKT[390]      = 144'hC4866D2061632074656D706F72206D657475;
        inPKT[391]      = 144'hC487732E205365642076656C207475727069;
        inPKT[392]      = 144'hC4887320666575676961742C20696163756C;
        inPKT[393]      = 144'hC489697320617567756520717569732C2074;
        inPKT[394]      = 144'hC48A696E636964756E74207475727069732E;
        inPKT[395]      = 144'hC48B0D0A0D0A566976616D757320706F7375;
        inPKT[396]      = 144'hC48C65726520706F72747469746F72206175;
        inPKT[397]      = 144'hC48D6775652C207661726975732061636375;
        inPKT[398]      = 144'hC48E6D73616E20656C69742076756C707574;
        inPKT[399]      = 144'hC48F61746520656765742E20517569737175;
        inPKT[400]      = 144'hC4906520736564206D616C65737561646120;
        inPKT[401]      = 144'hC4916E69736C2E20496E74657264756D2065;
        inPKT[402]      = 144'hC49274206D616C6573756164612066616D65;
        inPKT[403]      = 144'hC4937320616320616E746520697073756D20;
        inPKT[404]      = 144'hC4947072696D697320696E20666175636962;
        inPKT[405]      = 144'hC49575732E204E756E632074757270697320;
        inPKT[406]      = 144'hC4966469616D2C2073757363697069742061;
        inPKT[407]      = 144'hC497632065726F732076656C2C2074656D70;
        inPKT[408]      = 144'hC49875732076656E656E6174697320697073;
        inPKT[409]      = 144'hC499756D2E2044756973206C756374757320;
        inPKT[410]      = 144'hC49A72686F6E637573206D617373612E2046;
        inPKT[411]      = 144'hC49B75736365207574206C6163696E696120;
        inPKT[412]      = 144'hC49C7475727069732E20566976616D757320;
        inPKT[413]      = 144'hC49D72757472756D2074656C6C7573206175;
        inPKT[414]      = 144'hC49E6775652C206174206F726E617265206E;
        inPKT[415]      = 144'hC49F69736C20666163696C69736973206574;
        inPKT[416]      = 144'hC4A02E204E756E6320736564206E69736920;
        inPKT[417]      = 144'hC4A172697375732E20496E74656765722065;
        inPKT[418]      = 144'hC4A26C656D656E74756D206D617572697320;
        inPKT[419]      = 144'hC4A37175616D2C207574207665686963756C;
        inPKT[420]      = 144'hC4A461206D617572697320636F6E67756520;
        inPKT[421]      = 144'hC4A565752E0D0A0D0A467573636520612074;
        inPKT[422]      = 144'hC4A6656C6C75732073697420616D65742065;
        inPKT[423]      = 144'hC4A7726174206665726D656E74756D207363;
        inPKT[424]      = 144'hC4A8656C657269737175652E204375726162;
        inPKT[425]      = 144'hC4A96974757220696E2076656C6974206174;
        inPKT[426]      = 144'hC4AA20656E696D206C6163696E6961207665;
        inPKT[427]      = 144'hC4AB686963756C61206163206964206A7573;
        inPKT[428]      = 144'hC4AC746F2E2050726F696E206E6F6E20646F;
        inPKT[429]      = 144'hC4AD6C6F72206566666963697475722C2074;
        inPKT[430]      = 144'hC4AE696E636964756E74206F64696F206575;
        inPKT[431]      = 144'hC4AF2C20666175636962757320656E696D2E;
        inPKT[432]      = 144'hC4B02050656C6C656E746573717565206461;
        inPKT[433]      = 144'hC4B17069627573206F726369206163206C6F;
        inPKT[434]      = 144'hC4B272656D20696163756C69732C20736974;
        inPKT[435]      = 144'hC4B320616D657420626C616E646974206172;
        inPKT[436]      = 144'hC4B46375207472697374697175652E204165;
        inPKT[437]      = 144'hC4B56E65616E207472697374697175652074;
        inPKT[438]      = 144'hC4B66F72746F72206E6563206A7573746F20;
        inPKT[439]      = 144'hC4B7616C697175616D2C20696E2070726574;
        inPKT[440]      = 144'hC4B869756D2066656C6973206D6F6C657374;
        inPKT[441]      = 144'hC4B969652E205365642065742074656D7075;
        inPKT[442]      = 144'hC4BA732061756775652E204E756C6C612066;
        inPKT[443]      = 144'hC4BB72696E67696C6C6120656C656966656E;
        inPKT[444]      = 144'hC4BC6420697073756D207669766572726120;
        inPKT[445]      = 144'hC4BD6375727375732E20416C697175616D20;
        inPKT[446]      = 144'hC4BE6D6178696D7573206665726D656E7475;
        inPKT[447]      = 144'hC4BF6D206E69626820616320616363756D73;
        inPKT[448]      = 144'hC4C0616E2E204E756C6C6120666163696C69;
        inPKT[449]      = 144'hC4C173692E20566573746962756C756D2066;
        inPKT[450]      = 144'hC4C26163696C69736973206C656F20656765;
        inPKT[451]      = 144'hC4C3737461732073656D206D617474697320;
        inPKT[452]      = 144'hC4C4636F6E6775652E204D61757269732076;
        inPKT[453]      = 144'hC4C569746165206578206174207269737573;
        inPKT[454]      = 144'hC4C6206461706962757320656C656966656E;
        inPKT[455]      = 144'hC4C7642E20496E7465676572207574206572;
        inPKT[456]      = 144'hC4C86F7320636F6E6775652C20706F727474;
        inPKT[457]      = 144'hC4C969746F7220616E7465206E6F6E2C2069;
        inPKT[458]      = 144'hC4CA6E74657264756D20646F6C6F722E0D0A;
        inPKT[459]      = 144'hC4CB0D0A566573746962756C756D20656C65;
        inPKT[460]      = 144'hC4CC6966656E64206D617572697320657520;
        inPKT[461]      = 144'hC4CD6E6973692064696374756D2067726176;
        inPKT[462]      = 144'hC4CE6964612E2044756973206D6F6C6C6973;
        inPKT[463]      = 144'hC4CF206469616D2076656C20656E696D2074;
        inPKT[464]      = 144'hC4D0656D7075732C20766974616520646170;
        inPKT[465]      = 144'hC4D169627573206D61737361207361676974;
        inPKT[466]      = 144'hC4D27469732E204E756C6C61207574206175;
        inPKT[467]      = 144'hC4D363746F7220746F72746F722E204D6F72;
        inPKT[468]      = 144'hC4D4626920736564206C6F72656D2075726E;
        inPKT[469]      = 144'hC4D5612E204675736365206D61747469732C;
        inPKT[470]      = 144'hC4D6206D61676E6120616320636F6E64696D;
        inPKT[471]      = 144'hC4D7656E74756D20666575676961742C206D;
        inPKT[472]      = 144'hC4D86173736120647569206D6178696D7573;
        inPKT[473]      = 144'hC4D9206E756C6C612C20657520616C697175;
        inPKT[474]      = 144'hC4DA6574206E65717565206D617572697320;
        inPKT[475]      = 144'hC4DB6120657261742E205175697371756520;
        inPKT[476]      = 144'hC4DC617563746F722065737420757420696E;
        inPKT[477]      = 144'hC4DD74657264756D20636F6E736563746574;
        inPKT[478]      = 144'hC4DE75722E20446F6E656320656765742064;
        inPKT[479]      = 144'hC4DF69676E697373696D20746F72746F722C;
        inPKT[480]      = 144'hC4E02068656E647265726974206D61747469;
        inPKT[481]      = 144'hC4E17320657261742E2050656C6C656E7465;
        inPKT[482]      = 144'hC4E273717565206861626974616E74206D6F;
        inPKT[483]      = 144'hC4E372626920747269737469717565207365;
        inPKT[484]      = 144'hC4E46E6563747573206574206E6574757320;
        inPKT[485]      = 144'hC4E56574206D616C6573756164612066616D;
        inPKT[486]      = 144'hC4E665732061632074757270697320656765;
        inPKT[487]      = 144'hC4E7737461732E2051756973717565206F72;
        inPKT[488]      = 144'hC4E86E617265207661726975732074656D70;
        inPKT[489]      = 144'hC4E975732E0D0A0D0A4D6F72626920727574;
        inPKT[490]      = 144'hC4EA72756D20616E7465206E6962682C2061;
        inPKT[491]      = 144'hC4EB2076697665727261206E756C6C612068;
        inPKT[492]      = 144'hC4EC656E64726572697420696E2E2050726F;
        inPKT[493]      = 144'hC4ED696E2073757363697069742065676573;
        inPKT[494]      = 144'hC4EE74617320657261742C20757420617563;
        inPKT[495]      = 144'hC4EF746F72206F726369206D617474697320;
        inPKT[496]      = 144'hC4F0612E2050656C6C656E74657371756520;
        inPKT[497]      = 144'hC4F16C7563747573206672696E67696C6C61;
        inPKT[498]      = 144'hC4F220656C6974207574206C6163696E6961;
        inPKT[499]      = 144'hC4F32E205574206574206D61737361206E75;
        inPKT[500]      = 144'hC4F46C6C612E20536564206174206672696E;
        inPKT[501]      = 144'hC4F567696C6C61206C6F72656D2E2050726F;
        inPKT[502]      = 144'hC4F6696E206772617669646120616363756D;
        inPKT[503]      = 144'hC4F773616E20726973757320736564206269;
        inPKT[504]      = 144'hC4F862656E64756D2E204D616563656E6173;
        inPKT[505]      = 144'hC4F9206D616C657375616461206F64696F20;
        inPKT[506]      = 144'hC4FA75742076656C697420657569736D6F64;
        inPKT[507]      = 144'hC4FB20646170696275732E0D0A0D0A457469;
        inPKT[508]      = 144'hC4FC616D20636F6E677565206D6174746973;
        inPKT[509]      = 144'hC4FD20696163756C69732E204D6175726973;
        inPKT[510]      = 144'hC4FE20766974616520656666696369747572;
        inPKT[511]      = 144'hC4FF2073656D2E205365642070756C76696E;
        inPKT[512]      = 144'hC400617220646F6C6F72207574206D692065;
        inPKT[513]      = 144'hC4017569736D6F642068656E647265726974;
        inPKT[514]      = 144'hC4022E204E756C6C616D2061742067726176;
        inPKT[515]      = 144'hC40369646120646F6C6F722E204D6F726269;
        inPKT[516]      = 144'hC404206C656F207475727069732C20636F6E;
        inPKT[517]      = 144'hC405677565206E656320616C697175616D20;
        inPKT[518]      = 144'hC40675742C20636F6D6D6F646F20696E206E;
        inPKT[519]      = 144'hC407756E632E204E756C6C61206174206661;
        inPKT[520]      = 144'hC408756369627573206C656F2C2065752066;
        inPKT[521]      = 144'hC409657567696174206C616375732E204675;
        inPKT[522]      = 144'hC40A736365206E6F6E206567657374617320;
        inPKT[523]      = 144'hC40B7475727069732E205175697371756520;
        inPKT[524]      = 144'hC40C766974616520697073756D206D692E20;
        inPKT[525]      = 144'hC40D4E756E63206E6F6E206F726369207369;
        inPKT[526]      = 144'hC40E7420616D6574206E6973692076617269;
        inPKT[527]      = 144'hC40F757320706F72747469746F7220696E20;
        inPKT[528]      = 144'hC41076756C70757461746520746F72746F72;
        inPKT[529]      = 144'hC4112E204E756E6320636F6E76616C6C6973;
        inPKT[530]      = 144'hC4122067726176696461206469616D206120;
        inPKT[531]      = 144'hC413756C747269636965732E205175697371;
        inPKT[532]      = 144'hC4147565206575206A7573746F20636F6E64;
        inPKT[533]      = 144'hC415696D656E74756D2C2076617269757320;
        inPKT[534]      = 144'hC4166469616D2076656C2C20766573746962;
        inPKT[535]      = 144'hC417756C756D206D617373612E0D0A0D0A50;
        inPKT[536]      = 144'hC418656C6C656E7465737175652070656C6C;
        inPKT[537]      = 144'hC419656E7465737175652073617069656E20;
        inPKT[538]      = 144'hC41A6E657175652C20617563746F72206D61;
        inPKT[539]      = 144'hC41B6C65737561646120657261742068656E;
        inPKT[540]      = 144'hC41C647265726974206E65632E204E756C6C;
        inPKT[541]      = 144'hC41D6120706C616365726174206469616D20;
        inPKT[542]      = 144'hC41E68656E647265726974206D6173736120;
        inPKT[543]      = 144'hC41F626962656E64756D2C2061206D6F6C65;
        inPKT[544]      = 144'hC420737469652066656C69732068656E6472;
        inPKT[545]      = 144'hC421657269742E204D617572697320657569;
        inPKT[546]      = 144'hC422736D6F642076656E656E61746973206A;
        inPKT[547]      = 144'hC4237573746F2C20757420617563746F7220;
        inPKT[548]      = 144'hC424656C697420616C69717565742075742E;
        inPKT[549]      = 144'hC42520467573636520616C69717565742C20;
        inPKT[550]      = 144'hC4267175616D207574206469676E69737369;
        inPKT[551]      = 144'hC4276D2068656E6472657269742C206D6175;
        inPKT[552]      = 144'hC42872697320747572706973206469676E69;
        inPKT[553]      = 144'hC4297373696D20746F72746F722C20656765;
        inPKT[554]      = 144'hC42A742070656C6C656E7465737175652076;
        inPKT[555]      = 144'hC42B656C6974206F726369206E6563207175;
        inPKT[556]      = 144'hC42C616D2E204E756E632065676573746173;
        inPKT[557]      = 144'hC42D2070656C6C656E746573717565207269;
        inPKT[558]      = 144'hC42E7375732E204375726162697475722073;
        inPKT[559]      = 144'hC42F757363697069742074656D707573206C;
        inPKT[560]      = 144'hC430616375732C2065676574207072657469;
        inPKT[561]      = 144'hC431756D20656C69742074696E636964756E;
        inPKT[562]      = 144'hC43274206E6F6E2E20437261732075726E61;
        inPKT[563]      = 144'hC433206C6F72656D2C20706C616365726174;
        inPKT[564]      = 144'hC43420766F6C757470617420696D70657264;
        inPKT[565]      = 144'hC4356965742073697420616D65742C206567;
        inPKT[566]      = 144'hC43665737461732076656C206F7263692E0D;
        inPKT[567]      = 144'hC4370A0D0A50656C6C656E74657371756520;
        inPKT[568]      = 144'hC438736F64616C6573206665726D656E7475;
        inPKT[569]      = 144'hC4396D206E69736C2C206174206672696E67;
        inPKT[570]      = 144'hC43A696C6C61206475692073656D70657220;
        inPKT[571]      = 144'hC43B6665726D656E74756D2E204E756C6C61;
        inPKT[572]      = 144'hC43C6D20706C6163657261742076656C206D;
        inPKT[573]      = 144'hC43D692068656E64726572697420656C656D;
        inPKT[574]      = 144'hC43E656E74756D2E20457469616D206E6F6E;
        inPKT[575]      = 144'hC43F20697073756D2065782E204E616D2061;
        inPKT[576]      = 144'hC44063207363656C65726973717565206E69;
        inPKT[577]      = 144'hC44162682C2076656C20666163696C697369;
        inPKT[578]      = 144'hC44273206D692E20446F6E65632065676573;
        inPKT[579]      = 144'hC443746173206C616F726565742065726F73;
        inPKT[580]      = 144'hC4442C206567657420766F6C757470617420;
        inPKT[581]      = 144'hC4456D657475732E205072616573656E7420;
        inPKT[582]      = 144'hC446616363756D73616E20626962656E6475;
        inPKT[583]      = 144'hC4476D206E69736C206E65632076656E656E;
        inPKT[584]      = 144'hC448617469732E205365642072757472756D;
        inPKT[585]      = 144'hC449206D6920612073757363697069742070;
        inPKT[586]      = 144'hC44A686172657472612E2053656420736974;
        inPKT[587]      = 144'hC44B20616D657420696E74657264756D2074;
        inPKT[588]      = 144'hC44C75727069732E20416C697175616D2065;
        inPKT[589]      = 144'hC44D75206E69626820746F72746F722E2044;
        inPKT[590]      = 144'hC44E6F6E6563206661756369627573206461;
        inPKT[591]      = 144'hC44F7069627573206E6973692C2073656420;
        inPKT[592]      = 144'hC4506C616F72656574206F72636920736365;
        inPKT[593]      = 144'hC4516C6572697371756520696E2E0D0A0D0A;
        inPKT[594]      = 144'hC4524D617572697320696E2066656C697320;
        inPKT[595]      = 144'hC4536665726D656E74756D2C20636F6E7661;
        inPKT[596]      = 144'hC4546C6C69732061756775652076656C2C20;
        inPKT[597]      = 144'hC455706F7375657265206D692E2050656C6C;
        inPKT[598]      = 144'hC456656E746573717565207363656C657269;
        inPKT[599]      = 144'hC457737175652072686F6E637573206A7573;
        inPKT[600]      = 144'hC458746F2C2065752070756C76696E617220;
        inPKT[601]      = 144'hC459656E696D2070756C76696E6172207665;
        inPKT[602]      = 144'hC45A6C2E204D616563656E61732070686172;
        inPKT[603]      = 144'hC45B65747261206C696265726F206D61676E;
        inPKT[604]      = 144'hC45C612C20616320736F6C6C696369747564;
        inPKT[605]      = 144'hC45D696E206C656F206D6F6C6C6973206E6F;
        inPKT[606]      = 144'hC45E6E2E204E756C6C6120656C656D656E74;
        inPKT[607]      = 144'hC45F756D206F726E61726520656765737461;
        inPKT[608]      = 144'hC460732E20436C61737320617074656E7420;
        inPKT[609]      = 144'hC46174616369746920736F63696F73717520;
        inPKT[610]      = 144'hC4626164206C69746F726120746F72717565;
        inPKT[611]      = 144'hC4636E742070657220636F6E75626961206E;
        inPKT[612]      = 144'hC4646F737472612C2070657220696E636570;
        inPKT[613]      = 144'hC465746F732068696D656E61656F732E2050;
        inPKT[614]      = 144'hC46672616573656E74206175677565206D61;
        inPKT[615]      = 144'hC467757269732C2072686F6E637573207175;
        inPKT[616]      = 144'hC468697320657374206E6F6E2C206D6F6C6C;
        inPKT[617]      = 144'hC469697320636F6E76616C6C69732066656C;
        inPKT[618]      = 144'hC46A69732E2053757370656E646973736520;
        inPKT[619]      = 144'hC46B666163696C697369732C206F72636920;
        inPKT[620]      = 144'hC46C7669746165206C6163696E6961207465;
        inPKT[621]      = 144'hC46D6D706F722C206C656374757320736170;
        inPKT[622]      = 144'hC46E69656E206D6174746973207269737573;
        inPKT[623]      = 144'hC46F2C206E6F6E2073616769747469732065;
        inPKT[624]      = 144'hC4706C6974206E657175652071756973206A;
        inPKT[625]      = 144'hC4717573746F2E20446F6E6563206D616C65;
        inPKT[626]      = 144'hC4727375616461206C6163696E6961206475;
        inPKT[627]      = 144'hC473692E2050686173656C6C75732068656E;
        inPKT[628]      = 144'hC474647265726974206D6175726973206D61;
        inPKT[629]      = 144'hC475757269732C20736564206672696E6769;
        inPKT[630]      = 144'hC4766C6C61206C696265726F206672696E67;
        inPKT[631]      = 144'hC477696C6C6120696E2E2053656420617420;
        inPKT[632]      = 144'hC4786C6967756C6120696E206A7573746F20;
        inPKT[633]      = 144'hC47966696E696275732076756C7075746174;
        inPKT[634]      = 144'hC47A652E204E756E6320637572737573206E;
        inPKT[635]      = 144'hC47B657175652073697420616D6574206172;
        inPKT[636]      = 144'hC47C63752074696E636964756E742C207669;
        inPKT[637]      = 144'hC47D7461652070686172657472612073656D;
        inPKT[638]      = 144'hC47E20706F72747469746F722E20416C6971;
        inPKT[639]      = 144'hC47F75616D206D61747469732C206A757374;
        inPKT[640]      = 144'hC4806F206E6F6E20657569736D6F6420636F;
        inPKT[641]      = 144'hC4816E76616C6C69732C206E756E63206D69;
        inPKT[642]      = 144'hC48220636F6E736571756174206573742C20;
        inPKT[643]      = 144'hC4836E656320736F6C6C696369747564696E;
        inPKT[644]      = 144'hC484206C65637475732073617069656E2076;
        inPKT[645]      = 144'hC485656C206F64696F2E20496E2074656D70;
        inPKT[646]      = 144'hC4866F72206572617420646F6C6F722C2073;
        inPKT[647]      = 144'hC4876564207665686963756C612075726E61;
        inPKT[648]      = 144'hC48820636F6E736571756174207365642E0D;
        inPKT[649]      = 144'hC4890A0D0A4E616D2072686F6E6375732069;
        inPKT[650]      = 144'hC48A64206D6175726973206E656320646967;
        inPKT[651]      = 144'hC48B6E697373696D2E20496E20696D706572;
        inPKT[652]      = 144'hC48C6469657420756C747269636573206572;
        inPKT[653]      = 144'hC48D6174206E656320736F6C6C6963697475;
        inPKT[654]      = 144'hC48E64696E2E20496E746567657220736564;
        inPKT[655]      = 144'hC48F20636F6E64696D656E74756D2065726F;
        inPKT[656]      = 144'hC490732E20446F6E65632065676574206E75;
        inPKT[657]      = 144'hC4916E63206964206D617572697320747269;
        inPKT[658]      = 144'hC49273746971756520706F72747469746F72;
        inPKT[659]      = 144'hC493206C616F72656574207669746165206D;
        inPKT[660]      = 144'hC494657475732E204E756C6C612066616369;
        inPKT[661]      = 144'hC4956C6973692E204E756C6C616D20657520;
        inPKT[662]      = 144'hC4966C616375732061206469616D20747269;
        inPKT[663]      = 144'hC4977374697175652065676573746173206E;
        inPKT[664]      = 144'hC4986F6E20696163756C6973206D65747573;
        inPKT[665]      = 144'hC4992E20416C697175616D20696E2074656D;
        inPKT[666]      = 144'hC49A706F7220657261742C20696420636F6E;
        inPKT[667]      = 144'hC49B677565206D617373612E20566976616D;
        inPKT[668]      = 144'hC49C75732076656C20746F72746F72207669;
        inPKT[669]      = 144'hC49D746165206E69626820636F6D6D6F646F;
        inPKT[670]      = 144'hC49E206C6F626F7274697320717569732061;
        inPKT[671]      = 144'hC49F20697073756D2E2050726F696E20766F;
        inPKT[672]      = 144'hC4A06C7574706174207175616D206E6F6E20;
        inPKT[673]      = 144'hC4A166656C69732074656D7075732C206964;
        inPKT[674]      = 144'hC4A220706F737565726520646F6C6F722074;
        inPKT[675]      = 144'hC4A3656D706F722E205072616573656E7420;
        inPKT[676]      = 144'hC4A476697461652074696E636964756E7420;
        inPKT[677]      = 144'hC4A573617069656E2E204D616563656E6173;
        inPKT[678]      = 144'hC4A620666163696C69736973206D61747469;
        inPKT[679]      = 144'hC4A77320616E746520717569732076617269;
        inPKT[680]      = 144'hC4A875732E20446F6E65632070656C6C656E;
        inPKT[681]      = 144'hC4A97465737175652065726F732066657567;
        inPKT[682]      = 144'hC4AA6961742074696E636964756E7420636F;
        inPKT[683]      = 144'hC4AB6E64696D656E74756D2E2050726F696E;
        inPKT[684]      = 144'hC4AC20666175636962757320766F6C757470;
        inPKT[685]      = 144'hC4AD6174206D692073656420736167697474;
        inPKT[686]      = 144'hC4AE69732E0D0A0D0A447569732067726176;
        inPKT[687]      = 144'hC4AF69646120656C656D656E74756D20696E;
        inPKT[688]      = 144'hC4B074657264756D2E2050726F696E207369;
        inPKT[689]      = 144'hC4B17420616D6574207175616D206C696775;
        inPKT[690]      = 144'hC4B26C612E2050686173656C6C757320636F;
        inPKT[691]      = 144'hC4B36D6D6F646F2C2075726E6120696E2063;
        inPKT[692]      = 144'hC4B46F6E67756520766F6C75747061742C20;
        inPKT[693]      = 144'hC4B56C6967756C6120657820706861726574;
        inPKT[694]      = 144'hC4B67261206C6967756C612C20696E206469;
        inPKT[695]      = 144'hC4B76374756D206D61676E61206F72636920;
        inPKT[696]      = 144'hC4B86E6563206D61757269732E204E756E63;
        inPKT[697]      = 144'hC4B920617563746F7220636F6E7365637465;
        inPKT[698]      = 144'hC4BA74757220766F6C75747061742E204D6F;
        inPKT[699]      = 144'hC4BB7262692074696E636964756E74206E69;
        inPKT[700]      = 144'hC4BC626820757420656E696D206566666963;
        inPKT[701]      = 144'hC4BD6974757220677261766964612E204375;
        inPKT[702]      = 144'hC4BE72616269747572207669746165207175;
        inPKT[703]      = 144'hC4BF616D2065726F732E2044756973206672;
        inPKT[704]      = 144'hC4C0696E67696C6C6120616320746F72746F;
        inPKT[705]      = 144'hC4C17220696E2074696E636964756E742E20;
        inPKT[706]      = 144'hC4C24E756E632076656C206D617572697320;
        inPKT[707]      = 144'hC4C372697375732E20446F6E656320656C65;
        inPKT[708]      = 144'hC4C46966656E64206C6967756C6120736167;
        inPKT[709]      = 144'hC4C56974746973206E6973692066696E6962;
        inPKT[710]      = 144'hC4C675732C2061207363656C657269737175;
        inPKT[711]      = 144'hC4C765206C696265726F2070656C6C656E74;
        inPKT[712]      = 144'hC4C865737175652E20566573746962756C75;
        inPKT[713]      = 144'hC4C96D20747269737469717565206D617373;
        inPKT[714]      = 144'hC4CA61206E6962682C206174207665737469;
        inPKT[715]      = 144'hC4CB62756C756D206D61676E612066696E69;
        inPKT[716]      = 144'hC4CC6275732065752E0D0A0D0A4375726162;
        inPKT[717]      = 144'hC4CD6974757220696D706572646965742070;
        inPKT[718]      = 144'hC4CE757275732065676574206E756E632075;
        inPKT[719]      = 144'hC4CF6C7472696365732C2076697461652076;
        inPKT[720]      = 144'hC4D0656E656E61746973206D617373612063;
        inPKT[721]      = 144'hC4D16F6D6D6F646F2E2050656C6C656E7465;
        inPKT[722]      = 144'hC4D273717565206861626974616E74206D6F;
        inPKT[723]      = 144'hC4D372626920747269737469717565207365;
        inPKT[724]      = 144'hC4D46E6563747573206574206E6574757320;
        inPKT[725]      = 144'hC4D56574206D616C6573756164612066616D;
        inPKT[726]      = 144'hC4D665732061632074757270697320656765;
        inPKT[727]      = 144'hC4D7737461732E20496E206665726D656E74;
        inPKT[728]      = 144'hC4D8756D2061742075726E61206E6F6E2063;
        inPKT[729]      = 144'hC4D96F6E76616C6C69732E20446F6E656320;
        inPKT[730]      = 144'hC4DA6163206175677565206A7573746F2E20;
        inPKT[731]      = 144'hC4DB496E20617420656C6974206574206172;
        inPKT[732]      = 144'hC4DC6375206D6178696D7573206C75637475;
        inPKT[733]      = 144'hC4DD732E20467573636520657569736D6F64;
        inPKT[734]      = 144'hC4DE206E756E63206E65632076656E656E61;
        inPKT[735]      = 144'hC4DF74697320617563746F722E204C6F7265;
        inPKT[736]      = 144'hC4E06D20697073756D20646F6C6F72207369;
        inPKT[737]      = 144'hC4E17420616D65742C20636F6E7365637465;
        inPKT[738]      = 144'hC4E27475722061646970697363696E672065;
        inPKT[739]      = 144'hC4E36C69742E20446F6E6563206469637475;
        inPKT[740]      = 144'hC4E46D2074656D706F722072757472756D2E;
        inPKT[741]      = 144'hC4E52053656420656C656966656E64206469;
        inPKT[742]      = 144'hC4E6616D206964206D6173736120696D7065;
        inPKT[743]      = 144'hC4E772646965742C206163206F726E617265;
        inPKT[744]      = 144'hC4E8206C696265726F20656C656966656E64;
        inPKT[745]      = 144'hC4E92E204D616563656E6173206F726E6172;
        inPKT[746]      = 144'hC4EA65206D65747573206E756C6C612C2073;
        inPKT[747]      = 144'hC4EB697420616D6574206665726D656E7475;
        inPKT[748]      = 144'hC4EC6D20656C697420616C697175616D2069;
        inPKT[749]      = 144'hC4ED642E20446F6E656320756C7472696365;
        inPKT[750]      = 144'hC4EE7320746F72746F7220617420616E7465;
        inPKT[751]      = 144'hC4EF2068656E6472657269742C2065752073;
        inPKT[752]      = 144'hC4F061676974746973206A7573746F20756C;
        inPKT[753]      = 144'hC4F17472696365732E0D0A0D0A5072616573;
        inPKT[754]      = 144'hC4F2656E74206C7563747573207072657469;
        inPKT[755]      = 144'hC4F3756D206E657175652C2073697420616D;
        inPKT[756]      = 144'hC4F465742070656C6C656E74657371756520;
        inPKT[757]      = 144'hC4F56D617572697320656C656D656E74756D;
        inPKT[758]      = 144'hC4F6206E6F6E2E20557420626C616E646974;
        inPKT[759]      = 144'hC4F7207068617265747261206F64696F206E;
        inPKT[760]      = 144'hC4F86F6E20657569736D6F642E2051756973;
        inPKT[761]      = 144'hC4F9717565207669746165206C656F20616C;
        inPKT[762]      = 144'hC4FA697175616D2C20736F64616C65732074;
        inPKT[763]      = 144'hC4FB656C6C75732069642C20696163756C69;
        inPKT[764]      = 144'hC4FC73206D61757269732E204E616D206566;
        inPKT[765]      = 144'hC4FD6669636974757220696E207075727573;
        inPKT[766]      = 144'hC4FE2073656420616363756D73616E2E204D;
        inPKT[767]      = 144'hC4FF616563656E61732073697420616D6574;
        inPKT[768]      = 144'hC400206375727375732066656C69732E2051;
        inPKT[769]      = 144'hC4017569737175652066617563696275732C;
        inPKT[770]      = 144'hC4022064756920657420617563746F72206C;
        inPKT[771]      = 144'hC40375637475732C20616E74652065726174;
        inPKT[772]      = 144'hC40420706F73756572652065726F732C2075;
        inPKT[773]      = 144'hC4057420636F6E76616C6C6973206D657475;
        inPKT[774]      = 144'hC40673206C6563747573207669746165206C;
        inPKT[775]      = 144'hC407656F2E2053757370656E646973736520;
        inPKT[776]      = 144'hC408706F74656E74692E2043726173206574;
        inPKT[777]      = 144'hC40920646F6C6F72206E6F6E2075726E6120;
        inPKT[778]      = 144'hC40A7363656C657269737175652074726973;
        inPKT[779]      = 144'hC40B74697175652E20437261732072757472;
        inPKT[780]      = 144'hC40C756D206E65632076656C697420616320;
        inPKT[781]      = 144'hC40D73616769747469732E20446F6E656320;
        inPKT[782]      = 144'hC40E656C656966656E642C206C6163757320;
        inPKT[783]      = 144'hC40F7365642067726176696461206D616C65;
        inPKT[784]      = 144'hC41073756164612C20657820616E74652070;
        inPKT[785]      = 144'hC4116C616365726174206C65637475732C20;
        inPKT[786]      = 144'hC4126567657420636F6E677565206D617373;
        inPKT[787]      = 144'hC41361206D65747573206964206C61637573;
        inPKT[788]      = 144'hC4142E2053757370656E6469737365206964;
        inPKT[789]      = 144'hC4152072757472756D206C65637475732E20;
        inPKT[790]      = 144'hC4164675736365206D6178696D7573207365;
        inPKT[791]      = 144'hC41764206C6967756C612073656420766976;
        inPKT[792]      = 144'hC418657272612E204E616D206C7563747573;
        inPKT[793]      = 144'hC419206469616D20616E74652C2076697461;
        inPKT[794]      = 144'hC41A65206F726E617265206E657175652076;
        inPKT[795]      = 144'hC41B617269757320656765742E0D0A0D0A50;
        inPKT[796]      = 144'hC41C656C6C656E7465737175652061742065;
        inPKT[797]      = 144'hC41D6C6974206E6962682E20566573746962;
        inPKT[798]      = 144'hC41E756C756D20616E746520697073756D20;
        inPKT[799]      = 144'hC41F7072696D697320696E20666175636962;
        inPKT[800]      = 144'hC4207573206F726369206C75637475732065;
        inPKT[801]      = 144'hC4217420756C74726963657320706F737565;
        inPKT[802]      = 144'hC422726520637562696C6961204375726165;
        inPKT[803]      = 144'hC4233B204375726162697475722066617563;
        inPKT[804]      = 144'hC42469627573206469616D206C656F2C206E;
        inPKT[805]      = 144'hC425656320657569736D6F642073656D2065;
        inPKT[806]      = 144'hC42666666963697475722075742E20557420;
        inPKT[807]      = 144'hC4277665686963756C612061756775652061;
        inPKT[808]      = 144'hC42863206C696265726F20696163756C6973;
        inPKT[809]      = 144'hC4292C206E656320656C656966656E642065;
        inPKT[810]      = 144'hC42A7820706F7274612E204D6F7262692068;
        inPKT[811]      = 144'hC42B656E6472657269742067726176696461;
        inPKT[812]      = 144'hC42C2074696E636964756E742E2050726165;
        inPKT[813]      = 144'hC42D73656E7420646F6C6F72206C61637573;
        inPKT[814]      = 144'hC42E2C2074656D707573206575206672696E;
        inPKT[815]      = 144'hC42F67696C6C612073697420616D65742C20;
        inPKT[816]      = 144'hC430656C656966656E6420696E206E756C6C;
        inPKT[817]      = 144'hC431612E204E756C6C61206D6F6C6C697320;
        inPKT[818]      = 144'hC43265676574206D61676E61206E65632068;
        inPKT[819]      = 144'hC433656E6472657269742E20416C69717561;
        inPKT[820]      = 144'hC4346D20636F6E76616C6C69732073656D20;
        inPKT[821]      = 144'hC43576697461652073617069656E20646963;
        inPKT[822]      = 144'hC43674756D2C20757420766573746962756C;
        inPKT[823]      = 144'hC437756D206C6F72656D206672696E67696C;
        inPKT[824]      = 144'hC4386C612E20446F6E65632074656C6C7573;
        inPKT[825]      = 144'hC439206C696265726F2C2066657567696174;
        inPKT[826]      = 144'hC43A2075742066696E69627573206E65632C;
        inPKT[827]      = 144'hC43B20616C697175616D2073697420616D65;
        inPKT[828]      = 144'hC43C74206F7263692E204E756E6320737573;
        inPKT[829]      = 144'hC43D6369706974206E69736C206574206F72;
        inPKT[830]      = 144'hC43E6E61726520766573746962756C756D2E;
        inPKT[831]      = 144'hC43F204E756C6C616D206C6F626F72746973;
        inPKT[832]      = 144'hC4402073617069656E206A7573746F2C2073;
        inPKT[833]      = 144'hC441697420616D6574206469676E69737369;
        inPKT[834]      = 144'hC4426D206E756C6C6120636F6E64696D656E;
        inPKT[835]      = 144'hC44374756D20696E2E20536564206D6F6C65;
        inPKT[836]      = 144'hC4447374696520766F6C7574706174206E69;
        inPKT[837]      = 144'hC4457369206174206665726D656E74756D2E;
        inPKT[838]      = 144'hC446204E756C6C61206D6F6C657374696520;
        inPKT[839]      = 144'hC4476E697369207365642074757270697320;
        inPKT[840]      = 144'hC4486D6F6C65737469652C206E6F6E206961;
        inPKT[841]      = 144'hC44963756C6973206E756E63206661756369;
        inPKT[842]      = 144'hC44A6275732E2041656E65616E20696E7465;
        inPKT[843]      = 144'hC44B7264756D20706861726574726120636F;
        inPKT[844]      = 144'hC44C6E73656374657475722E20457469616D;
        inPKT[845]      = 144'hC44D206578206F7263692C20696163756C69;
        inPKT[846]      = 144'hC44E73206E6F6E20657569736D6F64206964;
        inPKT[847]      = 144'hC44F2C20756C6C616D636F72706572207363;
        inPKT[848]      = 144'hC450656C65726973717565206F64696F2E0D;
        inPKT[849]      = 144'hC4510A0D0A4E616D20756C74726963657320;
        inPKT[850]      = 144'hC452656C656966656E64206469616D2C2065;
        inPKT[851]      = 144'hC45367657420736F64616C65732073656D20;
        inPKT[852]      = 144'hC4546D61747469732061632E205574207665;
        inPKT[853]      = 144'hC4556E656E61746973206E69626820657520;
        inPKT[854]      = 144'hC4566C65637475732074696E636964756E74;
        inPKT[855]      = 144'hC4572064696374756D2E20566976616D7573;
        inPKT[856]      = 144'hC45820637572737573206175677565207175;
        inPKT[857]      = 144'hC4596973206C6F626F727469732065756973;
        inPKT[858]      = 144'hC45A6D6F642E204E756E6320616C69717561;
        inPKT[859]      = 144'hC45B6D206469616D20617420616E74652066;
        inPKT[860]      = 144'hC45C6163696C69736973206D6178696D7573;
        inPKT[861]      = 144'hC45D2E20457469616D20736564206C6F7265;
        inPKT[862]      = 144'hC45E6D206D61747469732C20636F6E76616C;
        inPKT[863]      = 144'hC45F6C69732075726E612076697461652C20;
        inPKT[864]      = 144'hC46074656D7075732073656D2E2056697661;
        inPKT[865]      = 144'hC4616D7573206567657374617320766F6C75;
        inPKT[866]      = 144'hC462747061742065726F7320657520756C74;
        inPKT[867]      = 144'hC46372696365732E20566573746962756C75;
        inPKT[868]      = 144'hC4646D20756C6C616D636F72706572206572;
        inPKT[869]      = 144'hC4656174206E756E632C206E6F6E2068656E;
        inPKT[870]      = 144'hC466647265726974206F64696F2070656C6C;
        inPKT[871]      = 144'hC467656E7465737175652069642E20467573;
        inPKT[872]      = 144'hC46863652075726E6120697073756D2C206C;
        inPKT[873]      = 144'hC4696163696E696120696E20737573636970;
        inPKT[874]      = 144'hC46A69742076656C2C2073656D7065722069;
        inPKT[875]      = 144'hC46B6E206F64696F2E2050656C6C656E7465;
        inPKT[876]      = 144'hC46C73717565206964206E696268206E6973;
        inPKT[877]      = 144'hC46D692E20416C697175616D20706F727461;
        inPKT[878]      = 144'hC46E206E69736C2065742065782069616375;
        inPKT[879]      = 144'hC46F6C6973207472697374697175652E2045;
        inPKT[880]      = 144'hC4707469616D206D61737361206F7263692C;
        inPKT[881]      = 144'hC471206567657374617320736564206C6F72;
        inPKT[882]      = 144'hC472656D20717569732C206469676E697373;
        inPKT[883]      = 144'hC473696D2073656D70657220616E74652E20;
        inPKT[884]      = 144'hC47453757370656E64697373652074696E63;
        inPKT[885]      = 144'hC4756964756E74206E6973692065782C2073;
        inPKT[886]      = 144'hC476656420766F6C75747061742065737420;
        inPKT[887]      = 144'hC4777661726975732076697461652E0D0A0D;
        inPKT[888]      = 144'hC4780A5365642073656D706572206C616369;
        inPKT[889]      = 144'hC4796E696120646F6C6F722E204E616D2075;
        inPKT[890]      = 144'hC47A742076656C697420696E206C61637573;
        inPKT[891]      = 144'hC47B20636F6E736563746574757220636F6E;
        inPKT[892]      = 144'hC47C76616C6C69732070656C6C656E746573;
        inPKT[893]      = 144'hC47D717565207365642073656D2E20537573;
        inPKT[894]      = 144'hC47E70656E646973736520636F6E64696D65;
        inPKT[895]      = 144'hC47F6E74756D20612065726F732069642075;
        inPKT[896]      = 144'hC4806C6C616D636F727065722E204D6F7262;
        inPKT[897]      = 144'hC48169206C75637475732075726E61207369;
        inPKT[898]      = 144'hC4827420616D657420657569736D6F642069;
        inPKT[899]      = 144'hC4836163756C69732E2050656C6C656E7465;
        inPKT[900]      = 144'hC4847371756520666163696C69736973206D;
        inPKT[901]      = 144'hC485617572697320657520656C656D656E74;
        inPKT[902]      = 144'hC486756D207661726975732E204F72636920;
        inPKT[903]      = 144'hC487766172697573206E61746F7175652070;
        inPKT[904]      = 144'hC488656E617469627573206574206D61676E;
        inPKT[905]      = 144'hC4896973206469732070617274757269656E;
        inPKT[906]      = 144'hC48A74206D6F6E7465732C206E6173636574;
        inPKT[907]      = 144'hC48B7572207269646963756C7573206D7573;
        inPKT[908]      = 144'hC48C2E20446F6E6563206469676E69737369;
        inPKT[909]      = 144'hC48D6D206120697073756D20756C74726963;
        inPKT[910]      = 144'hC48E6965732076656E656E617469732E2056;
        inPKT[911]      = 144'hC48F6976616D7573206E756E632076656C69;
        inPKT[912]      = 144'hC490742C207665686963756C612076697461;
        inPKT[913]      = 144'hC49165206D617373612075742C20636F6E76;
        inPKT[914]      = 144'hC492616C6C697320636F6E73656374657475;
        inPKT[915]      = 144'hC4937220746F72746F722E20517569737175;
        inPKT[916]      = 144'hC4946520616C697175616D2C206E69736C20;
        inPKT[917]      = 144'hC495636F6E67756520626C616E6469742075;
        inPKT[918]      = 144'hC4966C747269636965732C2075726E612074;
        inPKT[919]      = 144'hC4977572706973206D6174746973206D6167;
        inPKT[920]      = 144'hC4986E612C206E6F6E206665726D656E7475;
        inPKT[921]      = 144'hC4996D206475692076656C69742065752071;
        inPKT[922]      = 144'hC49A75616D2E0D0A0D0A496E207068617265;
        inPKT[923]      = 144'hC49B7472612076656C697420646F6C6F722C;
        inPKT[924]      = 144'hC49C20766974616520637572737573206F72;
        inPKT[925]      = 144'hC49D63692066696E696275732074696E6369;
        inPKT[926]      = 144'hC49E64756E742E20566976616D7573206964;
        inPKT[927]      = 144'hC49F20746F72746F722072686F6E6375732C;
        inPKT[928]      = 144'hC4A0207361676974746973206469616D2065;
        inPKT[929]      = 144'hC4A16765742C207072657469756D206D6175;
        inPKT[930]      = 144'hC4A27269732E2050686173656C6C75732065;
        inPKT[931]      = 144'hC4A36C656D656E74756D20656E696D206665;
        inPKT[932]      = 144'hC4A46C69732E204D6175726973206575206E;
        inPKT[933]      = 144'hC4A565717565206567657420707572757320;
        inPKT[934]      = 144'hC4A668656E64726572697420677261766964;
        inPKT[935]      = 144'hC4A7612E20416C697175616D206C69626572;
        inPKT[936]      = 144'hC4A86F206E6962682C20636F6E76616C6C69;
        inPKT[937]      = 144'hC4A9732061206E69736C2065742C2068656E;
        inPKT[938]      = 144'hC4AA64726572697420766573746962756C75;
        inPKT[939]      = 144'hC4AB6D2066656C69732E20446F6E65632065;
        inPKT[940]      = 144'hC4AC7569736D6F64206665726D656E74756D;
        inPKT[941]      = 144'hC4AD2074757270697320657520617563746F;
        inPKT[942]      = 144'hC4AE722E2041656E65616E20626962656E64;
        inPKT[943]      = 144'hC4AF756D2074757270697320696E206F6469;
        inPKT[944]      = 144'hC4B06F20636F6E76616C6C69732C20766974;
        inPKT[945]      = 144'hC4B1616520766172697573206578206C616F;
        inPKT[946]      = 144'hC4B2726565742E2046757363652076656C20;
        inPKT[947]      = 144'hC4B36D6920766974616520646F6C6F722066;
        inPKT[948]      = 144'hC4B46575676961742076756C707574617465;
        inPKT[949]      = 144'hC4B5206E6563207574206E756E632E204372;
        inPKT[950]      = 144'hC4B6617320646170696275732C20616E7465;
        inPKT[951]      = 144'hC4B7206964207665686963756C6120616C69;
        inPKT[952]      = 144'hC4B87175616D2C20656C69742065726F7320;
        inPKT[953]      = 144'hC4B97361676974746973206D692C206E6F6E;
        inPKT[954]      = 144'hC4BA20656C656966656E64206578206E756C;
        inPKT[955]      = 144'hC4BB6C6120656765742076656C69742E2053;
        inPKT[956]      = 144'hC4BC757370656E6469737365206964206469;
        inPKT[957]      = 144'hC4BD616D206475692E2053757370656E6469;
        inPKT[958]      = 144'hC4BE737365207072657469756D206A757374;
        inPKT[959]      = 144'hC4BF6F20736564206E69626820706F727474;
        inPKT[960]      = 144'hC4C069746F722C2076656C20696E74657264;
        inPKT[961]      = 144'hC4C1756D206D6175726973206D6178696D75;
        inPKT[962]      = 144'hC4C2732E20557420616C697175616D206C61;
        inPKT[963]      = 144'hC4C36375732070757275732C207369742061;
        inPKT[964]      = 144'hC4C46D657420696D70657264696574206E69;
        inPKT[965]      = 144'hC4C5626820666575676961742069642E2049;
        inPKT[966]      = 144'hC4C66E7465676572206C6F72656D206D6175;
        inPKT[967]      = 144'hC4C77269732C207072657469756D206E6F6E;
        inPKT[968]      = 144'hC4C8206E6973692065742C20646170696275;
        inPKT[969]      = 144'hC4C9732066696E69627573206F7263692E0D;
        inPKT[970]      = 144'hC4CA0A0D0A566573746962756C756D206961;
        inPKT[971]      = 144'hC4CB63756C69732C206D61676E6120617420;
        inPKT[972]      = 144'hC4CC6D6174746973206D6178696D75732C20;
        inPKT[973]      = 144'hC4CD61726375206572617420646170696275;
        inPKT[974]      = 144'hC4CE73206E756E632C206120766172697573;
        inPKT[975]      = 144'hC4CF206D657475732066656C697320736564;
        inPKT[976]      = 144'hC4D0206F7263692E204E756C6C616D206D69;
        inPKT[977]      = 144'hC4D1206E6962682C20656C656966656E6420;
        inPKT[978]      = 144'hC4D26E656320756C747269636573206E6563;
        inPKT[979]      = 144'hC4D32C20636F6E7365637465747572206163;
        inPKT[980]      = 144'hC4D420656E696D2E20536564206C75637475;
        inPKT[981]      = 144'hC4D5732073656D20717569732074656D706F;
        inPKT[982]      = 144'hC4D67220636F6E6775652E2053757370656E;
        inPKT[983]      = 144'hC4D7646973736520706F74656E74692E2045;
        inPKT[984]      = 144'hC4D87469616D2065676574206C696265726F;
        inPKT[985]      = 144'hC4D92076656C69742E204475697320766573;
        inPKT[986]      = 144'hC4DA746962756C756D20636F6E7365717561;
        inPKT[987]      = 144'hC4DB7420706F7274612E204D617572697320;
        inPKT[988]      = 144'hC4DC706F72747469746F7220747572706973;
        inPKT[989]      = 144'hC4DD20696E206D6173736120616C69717561;
        inPKT[990]      = 144'hC4DE6D20636F6E6775652E204E756C6C6120;
        inPKT[991]      = 144'hC4DF636F6E73656374657475722075726E61;
        inPKT[992]      = 144'hC4E0206D657475732C20696420696163756C;
        inPKT[993]      = 144'hC4E16973206E756E6320756C747269636965;
        inPKT[994]      = 144'hC4E27320656765742E204375726162697475;
        inPKT[995]      = 144'hC4E372206D6175726973206E657175652C20;
        inPKT[996]      = 144'hC4E4626962656E64756D207365642065726F;
        inPKT[997]      = 144'hC4E5732061742C206D6178696D757320756C;
        inPKT[998]      = 144'hC4E6747269636573207475727069732E0D0A;
        inPKT[999]      = 144'hC4E7496E74657264756D206574206D616C65;
        inPKT[1000]     = 144'hC4E873756164612066616D65732061632061;
        inPKT[1001]     = 144'hC4E96E746520697073756D207072696D6973;
        inPKT[1002]     = 144'hC4EA20696E2066617563696275732E205065;
        inPKT[1003]     = 144'hC4EB6C6C656E74657371756520736F6C6C69;
        inPKT[1004]     = 144'hC4EC6369747564696E20626C616E64697420;
        inPKT[1005]     = 144'hC4ED6665726D656E74756D2E2050656C6C65;
        inPKT[1006]     = 144'hC4EE6E746573717565206E6F6E206C696775;
        inPKT[1007]     = 144'hC4EF6C6120657520657261742076656E656E;
        inPKT[1008]     = 144'hC4F06174697320657569736D6F642E205065;
        inPKT[1009]     = 144'hC4F16C6C656E74657371756520736F64616C;
        inPKT[1010]     = 144'hC4F2657320766573746962756C756D20636F;
        inPKT[1011]     = 144'hC4F36E76616C6C69732E2050726F696E206D;
        inPKT[1012]     = 144'hC4F46F6C6573746965207072657469756D20;
        inPKT[1013]     = 144'hC4F565726F732076656C2065676573746173;
        inPKT[1014]     = 144'hC4F62E204D6F72626920736F6C6C69636974;
        inPKT[1015]     = 144'hC4F77564696E207075727573206163206665;
        inPKT[1016]     = 144'hC4F8726D656E74756D206D61747469732E20;
        inPKT[1017]     = 144'hC4F94E756E632076656C2074696E63696475;
        inPKT[1018]     = 144'hC4FA6E74206C696265726F2E204E756C6C61;
        inPKT[1019]     = 144'hC4FB20616C697175657420697073756D206E;
        inPKT[1020]     = 144'hC4FC6563207175616D20696D706572646965;
        inPKT[1021]     = 144'hC4FD7420696E74657264756D2E2050726165;
        inPKT[1022]     = 144'hC4FE73656E74206C6967756C612066656C69;
        inPKT[1023]     = 144'hC4FF732C20696163756C697320617420616C;
        inPKT[1024]     = 144'hC40069717565742061742C20736167697474;
        inPKT[1025]     = 144'hC4016973207175697320656C69742E0D0A51;
        inPKT[1026]     = 144'hC4027569737175652076656C20696D706572;
        inPKT[1027]     = 144'hC40364696574206E6962682E205068617365;
        inPKT[1028]     = 144'hC4046C6C75732072757472756D206469676E;
        inPKT[1029]     = 144'hC405697373696D207269737573206E6F6E20;
        inPKT[1030]     = 144'hC40674696E636964756E742E205665737469;
        inPKT[1031]     = 144'hC40762756C756D206E756E6320697073756D;
        inPKT[1032]     = 144'hC4082C2076656E656E617469732065676574;
        inPKT[1033]     = 144'hC40920706F72746120696E2C20636F6E7365;
        inPKT[1034]     = 144'hC40A63746574757220657520657261742E20;
        inPKT[1035]     = 144'hC40B446F6E6563207665686963756C612061;
        inPKT[1036]     = 144'hC40C6E74652076656C2072686F6E63757320;
        inPKT[1037]     = 144'hC40D66617563696275732E2050656C6C656E;
        inPKT[1038]     = 144'hC40E746573717565206A7573746F20746F72;
        inPKT[1039]     = 144'hC40F746F722C20766F6C757470617420696E;
        inPKT[1040]     = 144'hC410206D61757269732061742C2076617269;
        inPKT[1041]     = 144'hC41175732070686172657472612072697375;
        inPKT[1042]     = 144'hC412732E2051756973717565207574206469;
        inPKT[1043]     = 144'hC413616D2073757363697069742C20736F6C;
        inPKT[1044]     = 144'hC4146C696369747564696E2073617069656E;
        inPKT[1045]     = 144'hC4152065742C20696E74657264756D206C61;
        inPKT[1046]     = 144'hC4166375732E204D6F726269207269737573;
        inPKT[1047]     = 144'hC4172073656D2C2070656C6C656E74657371;
        inPKT[1048]     = 144'hC41875652065742074757270697320696E2C;
        inPKT[1049]     = 144'hC41920626C616E64697420736F6C6C696369;
        inPKT[1050]     = 144'hC41A747564696E2073656D2E205365642065;
        inPKT[1051]     = 144'hC41B6666696369747572206C696265726F20;
        inPKT[1052]     = 144'hC41C71756973207072657469756D20707265;
        inPKT[1053]     = 144'hC41D7469756D2E204E756C6C616D20617563;
        inPKT[1054]     = 144'hC41E746F72207361676974746973206C6F72;
        inPKT[1055]     = 144'hC41F656D2C20616320756C74726963657320;
        inPKT[1056]     = 144'hC42061726375206D6178696D757320656765;
        inPKT[1057]     = 144'hC421742E0D0A566573746962756C756D2076;
        inPKT[1058]     = 144'hC4226F6C7574706174206C6967756C612061;
        inPKT[1059]     = 144'hC4237563746F722073656D20766976657272;
        inPKT[1060]     = 144'hC424612C20756C6C616D636F727065722065;
        inPKT[1061]     = 144'hC4257569736D6F64206E6571756520706F72;
        inPKT[1062]     = 144'hC426747469746F722E2053757370656E6469;
        inPKT[1063]     = 144'hC4277373652076697665727261207363656C;
        inPKT[1064]     = 144'hC42865726973717565206F64696F2072686F;
        inPKT[1065]     = 144'hC4296E63757320766F6C75747061742E2041;
        inPKT[1066]     = 144'hC42A6C697175616D206572617420766F6C75;
        inPKT[1067]     = 144'hC42B747061742E2053757370656E64697373;
        inPKT[1068]     = 144'hC42C6520706F74656E74692E20496E206861;
        inPKT[1069]     = 144'hC42D632068616269746173736520706C6174;
        inPKT[1070]     = 144'hC42E65612064696374756D73742E2050726F;
        inPKT[1071]     = 144'hC42F696E207574206E756C6C612075742064;
        inPKT[1072]     = 144'hC4307569207363656C657269737175652064;
        inPKT[1073]     = 144'hC431696374756D2E20517569737175652073;
        inPKT[1074]     = 144'hC43275736369706974206E69626820706F73;
        inPKT[1075]     = 144'hC43375657265207175616D2076756C707574;
        inPKT[1076]     = 144'hC4346174652C206575206C6163696E696120;
        inPKT[1077]     = 144'hC435616E746520677261766964612E204375;
        inPKT[1078]     = 144'hC43672616269747572206D61737361206C6F;
        inPKT[1079]     = 144'hC43772656D2C206F726E617265206575206D;
        inPKT[1080]     = 144'hC4386F6C6C69732061742C20706861726574;
        inPKT[1081]     = 144'hC4397261206E6563206D617373612E204E75;
        inPKT[1082]     = 144'hC43A6C6C612066696E6962757320656C6569;
        inPKT[1083]     = 144'hC43B66656E64206F7263692073697420616D;
        inPKT[1084]     = 144'hC43C657420636F6E73656374657475722E20;
        inPKT[1085]     = 144'hC43D5365642074656D707573207669746165;
        inPKT[1086]     = 144'hC43E2061726375206E6563206665726D656E;
        inPKT[1087]     = 144'hC43F74756D2E2041656E65616E2070656C6C;
        inPKT[1088]     = 144'hC440656E7465737175652076697461652064;
        inPKT[1089]     = 144'hC4416F6C6F7220696E20616363756D73616E;
        inPKT[1090]     = 144'hC4422E2043726173206469676E697373696D;
        inPKT[1091]     = 144'hC4432076756C707574617465206D6F6C6C69;
        inPKT[1092]     = 144'hC444732E204D617572697320706F72746120;
        inPKT[1093]     = 144'hC44576656E656E617469732072697375732C;
        inPKT[1094]     = 144'hC4462065752074726973746971756520646F;
        inPKT[1095]     = 144'hC4476C6F722072757472756D20696E2E2046;
        inPKT[1096]     = 144'hC4487573636520636F6E64696D656E74756D;
        inPKT[1097]     = 144'hC449206F7263692066656C69732C20736974;
        inPKT[1098]     = 144'hC44A20616D657420636F6E76616C6C697320;
        inPKT[1099]     = 144'hC44B6C696265726F2074696E636964756E74;
        inPKT[1100]     = 144'hC44C2061632E0D0A566573746962756C756D;
        inPKT[1101]     = 144'hC44D20696D7065726469657420656C697420;
        inPKT[1102]     = 144'hC44E74656D706F72207175616D2067726176;
        inPKT[1103]     = 144'hC44F6964612C207574206D616C6573756164;
        inPKT[1104]     = 144'hC450612074656C6C757320696D7065726469;
        inPKT[1105]     = 144'hC45165742E2050686173656C6C7573206F64;
        inPKT[1106]     = 144'hC452696F2073656D2C206D61747469732073;
        inPKT[1107]     = 144'hC453656420756C7472696365732061742C20;
        inPKT[1108]     = 144'hC454766976657272612076656C206475692E;
        inPKT[1109]     = 144'hC455204E756E632075726E61206D65747573;
        inPKT[1110]     = 144'hC4562C206C7563747573206163206D617869;
        inPKT[1111]     = 144'hC4576D757320696E2C20636F6E7365637465;
        inPKT[1112]     = 144'hC458747572206E6F6E206E6973692E204E75;
        inPKT[1113]     = 144'hC4596C6C612073697420616D657420626962;
        inPKT[1114]     = 144'hC45A656E64756D2076656C69742E20446F6E;
        inPKT[1115]     = 144'hC45B6563207175697320656E696D206E6F6E;
        inPKT[1116]     = 144'hC45C20726973757320626C616E6469742066;
        inPKT[1117]     = 144'hC45D6163696C697369732071756973206E65;
        inPKT[1118]     = 144'hC45E632072697375732E2043757261626974;
        inPKT[1119]     = 144'hC45F75722065752065737420766974616520;
        inPKT[1120]     = 144'hC4606C656374757320626C616E6469742061;
        inPKT[1121]     = 144'hC4616C69717565742E20566573746962756C;
        inPKT[1122]     = 144'hC462756D20616E746520697073756D207072;
        inPKT[1123]     = 144'hC463696D697320696E206661756369627573;
        inPKT[1124]     = 144'hC464206F726369206C756374757320657420;
        inPKT[1125]     = 144'hC465756C74726963657320706F7375657265;
        inPKT[1126]     = 144'hC46620637562696C69612043757261653B20;
        inPKT[1127]     = 144'hC467566573746962756C756D206163206469;
        inPKT[1128]     = 144'hC468676E697373696D206E756E632E205175;
        inPKT[1129]     = 144'hC469697371756520696E2073616769747469;
        inPKT[1130]     = 144'hC46A732074656C6C75732C2073697420616D;
        inPKT[1131]     = 144'hC46B6574206665726D656E74756D206E6962;
        inPKT[1132]     = 144'hC46C682E0D0A496E206469676E697373696D;
        inPKT[1133]     = 144'hC46D20726973757320766974616520707572;
        inPKT[1134]     = 144'hC46E757320766573746962756C756D2C2061;
        inPKT[1135]     = 144'hC46F7420656C656D656E74756D206E756C6C;
        inPKT[1136]     = 144'hC4706120706F73756572652E20536564206D;
        inPKT[1137]     = 144'hC4716174746973206E756E63206E6962682E;
        inPKT[1138]     = 144'hC4722053757370656E64697373652070656C;
        inPKT[1139]     = 144'hC4736C656E74657371756520706C61636572;
        inPKT[1140]     = 144'hC4746174207363656C657269737175652E20;
        inPKT[1141]     = 144'hC47541656E65616E2066657567696174206D;
        inPKT[1142]     = 144'hC476617572697320696420636F6E67756520;
        inPKT[1143]     = 144'hC4776C6163696E69612E20457469616D2073;
        inPKT[1144]     = 144'hC47875736369706974206C6967756C612074;
        inPKT[1145]     = 144'hC479656C6C75732C206120636F6E67756520;
        inPKT[1146]     = 144'hC47A6C656374757320616C697175616D2076;
        inPKT[1147]     = 144'hC47B65686963756C612E2053757370656E64;
        inPKT[1148]     = 144'hC47C69737365206567657420616E74652076;
        inPKT[1149]     = 144'hC47D656C20656E696D206D616C6573756164;
        inPKT[1150]     = 144'hC47E6120766976657272612E2050726F696E;
        inPKT[1151]     = 144'hC47F2074696E636964756E74206172637520;
        inPKT[1152]     = 144'hC480656765742076756C7075746174652061;
        inPKT[1153]     = 144'hC4816363756D73616E2E20496E2076697461;
        inPKT[1154]     = 144'hC48265206469616D206E6962682E204D6F72;
        inPKT[1155]     = 144'hC4836269206D6178696D75732066656C6973;
        inPKT[1156]     = 144'hC48420696420636F6E736563746574757220;
        inPKT[1157]     = 144'hC485616C697175616D2E204E756C6C612066;
        inPKT[1158]     = 144'hC4866163696C6973692E0D0A566573746962;
        inPKT[1159]     = 144'hC487756C756D20766573746962756C756D20;
        inPKT[1160]     = 144'hC48865666669636974757220746F72746F72;
        inPKT[1161]     = 144'hC4892073697420616D657420666163696C69;
        inPKT[1162]     = 144'hC48A7369732E204D616563656E6173206E6F;
        inPKT[1163]     = 144'hC48B6E2074656C6C7573206F7263692E2050;
        inPKT[1164]     = 144'hC48C686173656C6C7573206E6F6E206C7563;
        inPKT[1165]     = 144'hC48D747573206A7573746F2C206174207375;
        inPKT[1166]     = 144'hC48E7363697069742074656C6C75732E2046;
        inPKT[1167]     = 144'hC48F757363652068656E647265726974206E;
        inPKT[1168]     = 144'hC4906563206E6962682076656C2063757273;
        inPKT[1169]     = 144'hC49175732E2053757370656E646973736520;
        inPKT[1170]     = 144'hC492706F74656E74692E2044756973206C69;
        inPKT[1171]     = 144'hC49367756C612066656C69732C2065666669;
        inPKT[1172]     = 144'hC49463697475722065742076656C69742061;
        inPKT[1173]     = 144'hC495742C20666163696C6973697320636F6E;
        inPKT[1174]     = 144'hC49676616C6C6973206A7573746F2E204E75;
        inPKT[1175]     = 144'hC4976C6C616D206C6F626F72746973207065;
        inPKT[1176]     = 144'hC4986C6C656E74657371756520736F6C6C69;
        inPKT[1177]     = 144'hC4996369747564696E2E204E616D20736974;
        inPKT[1178]     = 144'hC49A20616D657420646F6C6F722073697420;
        inPKT[1179]     = 144'hC49B616D6574206C656374757320696D7065;
        inPKT[1180]     = 144'hC49C726469657420636F6E7365717561742E;
        inPKT[1181]     = 144'hC49D20416C697175616D206C756374757320;
        inPKT[1182]     = 144'hC49E7363656C657269737175652070757275;
        inPKT[1183]     = 144'hC49F732C206964206672696E67696C6C6120;
        inPKT[1184]     = 144'hC4A073656D20766F6C75747061742061632E;
        inPKT[1185]     = 144'hC4A1205365642074656D706F722C20656E69;
        inPKT[1186]     = 144'hC4A26D206567657420657569736D6F642066;
        inPKT[1187]     = 144'hC4A36163696C697369732C206E6973692065;
        inPKT[1188]     = 144'hC4A4782073656D70657220697073756D2C20;
        inPKT[1189]     = 144'hC4A5696E207361676974746973206F726369;
        inPKT[1190]     = 144'hC4A6207175616D20696E206C65637475732E;
        inPKT[1191]     = 144'hC4A720557420766974616520656C6974206C;
        inPKT[1192]     = 144'hC4A86967756C612E204E756E632065676573;
        inPKT[1193]     = 144'hC4A97461732C206D69207669746165206961;
        inPKT[1194]     = 144'hC4AA63756C6973206D61747469732C206475;
        inPKT[1195]     = 144'hC4AB69206E69626820656C656966656E6420;
        inPKT[1196]     = 144'hC4AC6E69736C2C206567657420706F727461;
        inPKT[1197]     = 144'hC4AD206C696265726F206175677565207175;
        inPKT[1198]     = 144'hC4AE697320656E696D2E2053656420736974;
        inPKT[1199]     = 144'hC4AF20616D65742070756C76696E61722065;
        inPKT[1200]     = 144'hC4B0782C2076656C2070656C6C656E746573;
        inPKT[1201]     = 144'hC4B1717565206C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
