`include "SIMON_defintions.svh"

module test_SIMON_128128_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 600
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 272'hE7000F0E0D0C0B0A0908070605040302010000000000000000000000000000000000;
        inPKT[1]        = 272'hC7014C6F72656D20697073756D20646F6C6F722073697420616D65742C20636F6E73;
        inPKT[2]        = 272'hC702656374657475722061646970697363696E6720656C69742E2043757261626974;
        inPKT[3]        = 272'hC703757220756C6C616D636F727065722074656D707573206E6973692C2065742070;
        inPKT[4]        = 272'hC7046F73756572652075726E612E2041656E65616E20736564206772617669646120;
        inPKT[5]        = 272'hC7056C616375732E204E756C6C6120666163696C6973692E204E756C6C612074656D;
        inPKT[6]        = 272'hC706707573206F726369207175697320656C697420666575676961742C2076656C20;
        inPKT[7]        = 272'hC70773656D706572206C656F20696D706572646965742E204D616563656E61732065;
        inPKT[8]        = 272'hC70874206E756E6320696E206E69626820666163696C6973697320636F6E76616C6C;
        inPKT[9]        = 272'hC70969732E2053656420636F6E6775652068656E64726572697420696163756C6973;
        inPKT[10]       = 272'hC70A2E20566976616D7573207665686963756C61206C7563747573206573742C2076;
        inPKT[11]       = 272'hC70B69746165207375736369706974206E69736C20706F72747469746F722061632E;
        inPKT[12]       = 272'hC70C0D0A0D0A446F6E6563206D6F6C65737469652073617069656E2069642076756C;
        inPKT[13]       = 272'hC70D70757461746520766573746962756C756D2E204E756C6C6120696E206C696775;
        inPKT[14]       = 272'hC70E6C61206672696E67696C6C612C20756C6C616D636F727065722075726E612065;
        inPKT[15]       = 272'hC70F742C20706F72747469746F72206C65637475732E205175697371756520626C61;
        inPKT[16]       = 272'hC7106E646974206575206D61757269732061632068656E6472657269742E204E756C;
        inPKT[17]       = 272'hC7116C612076656E656E617469732C206D65747573206574206C7563747573206672;
        inPKT[18]       = 272'hC712696E67696C6C612C206E6962682076656C697420756C6C616D636F7270657220;
        inPKT[19]       = 272'hC7136469616D2C20656765742065666669636974757220697073756D207475727069;
        inPKT[20]       = 272'hC71473206174206E6962682E2055742065676574207072657469756D2065726F732C;
        inPKT[21]       = 272'hC71520656765742064696374756D206C616375732E204D616563656E617320757420;
        inPKT[22]       = 272'hC716656E696D2065782E2041656E65616E2076697461652073656D7065722066656C;
        inPKT[23]       = 272'hC71769732C2073656420756C747269636965732072697375732E20446F6E65632063;
        inPKT[24]       = 272'hC7186F6E7365637465747572206D69206E69736C2C20617420637572737573206970;
        inPKT[25]       = 272'hC71973756D206772617669646120612E2050686173656C6C75732073697420616D65;
        inPKT[26]       = 272'hC71A74206D61676E612076656C20697073756D206567657374617320706F7274612E;
        inPKT[27]       = 272'hC71B20566976616D7573206C756374757320656E696D20656765742074656D706F72;
        inPKT[28]       = 272'hC71C2073616769747469732E20416C697175616D20626962656E64756D2073656D20;
        inPKT[29]       = 272'hC71D6120636F6E7365637465747572206566666963697475722E20446F6E65632073;
        inPKT[30]       = 272'hC71E63656C6572697371756520616C697175616D206375727375732E204375726162;
        inPKT[31]       = 272'hC71F697475722073697420616D657420626962656E64756D20656C69742E20536564;
        inPKT[32]       = 272'hC720206469616D206A7573746F2C20696163756C69732071756973206E756C6C6120;
        inPKT[33]       = 272'hC72176697461652C20616C697175616D20657569736D6F642066656C69732E0D0A0D;
        inPKT[34]       = 272'hC7220A50726F696E20646170696275732C206469616D2076756C7075746174652066;
        inPKT[35]       = 272'hC72372696E67696C6C61206D616C6573756164612C206A7573746F20707572757320;
        inPKT[36]       = 272'hC724636F6D6D6F646F20646F6C6F722C2075742064696374756D2065726174206E75;
        inPKT[37]       = 272'hC7256E632072757472756D2075726E612E204E756C6C612067726176696461207572;
        inPKT[38]       = 272'hC7266E6120766974616520696D70657264696574206C616F726565742E2050656C6C;
        inPKT[39]       = 272'hC727656E7465737175652072686F6E63757320626962656E64756D206E6962682C20;
        inPKT[40]       = 272'hC7286964206D6F6C6C6973206469616D2073757363697069742061632E2050656C6C;
        inPKT[41]       = 272'hC729656E7465737175652076656C20696163756C6973206475692E204D6F72626920;
        inPKT[42]       = 272'hC72A617420616C6971756574206D617373612E2050726F696E207669746165206F72;
        inPKT[43]       = 272'hC72B6E617265206F64696F2C2065752076756C70757461746520697073756D2E2050;
        inPKT[44]       = 272'hC72C726F696E206C6F626F727469732C2073656D206E656320657569736D6F642074;
        inPKT[45]       = 272'hC72D696E636964756E742C206175677565206D6175726973207363656C6572697371;
        inPKT[46]       = 272'hC72E7565206D61676E612C20657420706F7375657265206D69206E69736C206E6563;
        inPKT[47]       = 272'hC72F206E6973692E20467573636520656C6974206E657175652C2076617269757320;
        inPKT[48]       = 272'hC7306574206672696E67696C6C612076697461652C207661726975732076656C206E;
        inPKT[49]       = 272'hC731657175652E204E756C6C612065742074656D707573206A7573746F2E204D6F72;
        inPKT[50]       = 272'hC732626920756C6C616D636F7270657220737573636970697420636F6E6775652E20;
        inPKT[51]       = 272'hC73353656420656C656966656E64206F64696F206163207375736369706974206469;
        inPKT[52]       = 272'hC734676E697373696D2E205175697371756520616E746520656E696D2C20626C616E;
        inPKT[53]       = 272'hC73564697420696E20636F6E7365717561742061632C20696E74657264756D207669;
        inPKT[54]       = 272'hC7367461652070757275732E204D617572697320657569736D6F6420706F73756572;
        inPKT[55]       = 272'hC73765206C65637475732E20566976616D757320696E74657264756D207175616D20;
        inPKT[56]       = 272'hC73865752073656D7065722066617563696275732E0D0A0D0A496E206D6F6C657374;
        inPKT[57]       = 272'hC7396965206E756C6C6120616E74652C20616320696E74657264756D206D61676E61;
        inPKT[58]       = 272'hC73A20636F6E64696D656E74756D20636F6E64696D656E74756D2E20447569732075;
        inPKT[59]       = 272'hC73B6C7472696369657320736F64616C6573206E756C6C612C2073697420616D6574;
        inPKT[60]       = 272'hC73C20756C6C616D636F72706572206F64696F207072657469756D206E65632E2046;
        inPKT[61]       = 272'hC73D75736365207365642072697375732070656C6C656E7465737175652C20636F6E;
        inPKT[62]       = 272'hC73E76616C6C69732073656D20656765742C2068656E64726572697420657261742E;
        inPKT[63]       = 272'hC73F204D6F72626920736F64616C6573207665686963756C61206C6F626F72746973;
        inPKT[64]       = 272'hC7402E2041656E65616E206120746F72746F72206375727375732C207363656C6572;
        inPKT[65]       = 272'hC7416973717565206C6967756C6120706F72747469746F722C206567657374617320;
        inPKT[66]       = 272'hC74265726F732E20447569732074696E636964756E7420746F72746F722069642070;
        inPKT[67]       = 272'hC7436F737565726520677261766964612E20496E20636F6E76616C6C6973206D6920;
        inPKT[68]       = 272'hC744696420697073756D206D616C6573756164612C2075742064696374756D206572;
        inPKT[69]       = 272'hC7456F7320696D706572646965742E2050726F696E20756C6C616D636F727065722C;
        inPKT[70]       = 272'hC746206D61757269732069642076617269757320636F6E6775652C2065726F732073;
        inPKT[71]       = 272'hC747617069656E2072686F6E637573206D692C20617420617563746F72206E657175;
        inPKT[72]       = 272'hC748652061726375206C616F72656574206469616D2E0D0A0D0A467573636520706F;
        inPKT[73]       = 272'hC74972747469746F72206C696265726F20617263752C206C6163696E69612068656E;
        inPKT[74]       = 272'hC74A647265726974206469616D20636F6E76616C6C6973207365642E205068617365;
        inPKT[75]       = 272'hC74B6C6C7573206E6F6E207475727069732070686172657472612C20756C6C616D63;
        inPKT[76]       = 272'hC74C6F72706572206E657175652076656C2C20736F6C6C696369747564696E207665;
        inPKT[77]       = 272'hC74D6C69742E2050656C6C656E746573717565206861626974616E74206D6F726269;
        inPKT[78]       = 272'hC74E207472697374697175652073656E6563747573206574206E6574757320657420;
        inPKT[79]       = 272'hC74F6D616C6573756164612066616D65732061632074757270697320656765737461;
        inPKT[80]       = 272'hC750732E204E616D206E65632073617069656E206D6F6C65737469652C2064696374;
        inPKT[81]       = 272'hC751756D206D6173736120656765742C2065676573746173206F64696F2E20457469;
        inPKT[82]       = 272'hC752616D20617263752073617069656E2C207072657469756D2061206D6F6C6C6973;
        inPKT[83]       = 272'hC75320612C2076756C707574617465206E6F6E20657261742E205574207669746165;
        inPKT[84]       = 272'hC754206E696268206C6F626F72746973206C65637475732066617563696275732070;
        inPKT[85]       = 272'hC7556F7274612065752073697420616D6574206E69736C2E204D6F72626920706F72;
        inPKT[86]       = 272'hC756747469746F722076656C697420657520646F6C6F72206C616F726565742C2073;
        inPKT[87]       = 272'hC757697420616D657420696D7065726469657420656E696D20736F64616C65732E20;
        inPKT[88]       = 272'hC7584E756C6C616D20756C6C616D636F72706572207475727069732061742070656C;
        inPKT[89]       = 272'hC7596C656E746573717565207661726975732E20566976616D757320657520696D70;
        inPKT[90]       = 272'hC75A657264696574206E657175652E20536564207175697320617563746F7220616E;
        inPKT[91]       = 272'hC75B74652E204D61757269732073656D70657220697073756D207365642064756920;
        inPKT[92]       = 272'hC75C706F73756572652C20617420616C697175616D206D6574757320656C65696665;
        inPKT[93]       = 272'hC75D6E642E204E756C6C616D2074726973746971756520656C656966656E64206572;
        inPKT[94]       = 272'hC75E6F732C2065676574206665726D656E74756D20697073756D20656C656D656E74;
        inPKT[95]       = 272'hC75F756D206E65632E0D0A0D0A50656C6C656E7465737175652068656E6472657269;
        inPKT[96]       = 272'hC7607420626962656E64756D206C6967756C612C20657420736F64616C6573206D61;
        inPKT[97]       = 272'hC761676E61206461706962757320696E2E20496E20616C697175657420746F72746F;
        inPKT[98]       = 272'hC76272206567657420636F6E736563746574757220636F6E73656374657475722E20;
        inPKT[99]       = 272'hC763517569737175652074726973746971756520726973757320657261742C206574;
        inPKT[100]      = 272'hC76420616C697175657420656C697420616C69717565742065752E20496E74656765;
        inPKT[101]      = 272'hC76572206E6F6E206D61676E6120696E2066656C697320706F72747469746F722073;
        inPKT[102]      = 272'hC766616769747469732E20517569737175652076697665727261206F726369206163;
        inPKT[103]      = 272'hC7672072757472756D206C616F726565742E2041656E65616E20636F6E76616C6C69;
        inPKT[104]      = 272'hC768732064696374756D207475727069732C2065742066696E696275732073617069;
        inPKT[105]      = 272'hC769656E20636F6E67756520696E2E2053656420612065726174206F726E6172652C;
        inPKT[106]      = 272'hC76A206D6F6C6C6973206E69736C2061632C206469676E697373696D206E65717565;
        inPKT[107]      = 272'hC76B2E2051756973717565206D616C65737561646120706F73756572652074757270;
        inPKT[108]      = 272'hC76C697320657520756C6C616D636F727065722E20446F6E65632076697665727261;
        inPKT[109]      = 272'hC76D20626962656E64756D206E756E632C2064696374756D20696D70657264696574;
        inPKT[110]      = 272'hC76E206E65717565206D6178696D757320696E2E20446F6E656320757420756C7472;
        inPKT[111]      = 272'hC76F6963657320646F6C6F722E20566976616D757320736564206175677565207072;
        inPKT[112]      = 272'hC770657469756D2C20766F6C757470617420657261742061632C20706F7274612064;
        inPKT[113]      = 272'hC77169616D2E204D617572697320696E20707572757320756C747269636965732C20;
        inPKT[114]      = 272'hC7727375736369706974206469616D207365642C2074696E636964756E7420656E69;
        inPKT[115]      = 272'hC7736D2E20446F6E6563207175697320706F7375657265206E6962682E20496E2068;
        inPKT[116]      = 272'hC77461632068616269746173736520706C617465612064696374756D73742E0D0A0D;
        inPKT[117]      = 272'hC7750A4D6F726269206F726E617265206A7573746F206174207175616D2066617563;
        inPKT[118]      = 272'hC776696275732C2073697420616D6574206D6F6C6573746965206C656F2063757273;
        inPKT[119]      = 272'hC77775732E204D6175726973206C616F7265657420616E74652061206D6574757320;
        inPKT[120]      = 272'hC778656666696369747572207661726975732E205365642076656C206F7263692073;
        inPKT[121]      = 272'hC77961676974746973206E756E6320626C616E64697420636F6E7365717561742E20;
        inPKT[122]      = 272'hC77A5072616573656E74206D616C657375616461206E657175652071756973206469;
        inPKT[123]      = 272'hC77B6374756D206469676E697373696D2E20446F6E656320666163696C6973697320;
        inPKT[124]      = 272'hC77C73697420616D65742076656C6974206575206C6F626F727469732E204E756C6C;
        inPKT[125]      = 272'hC77D616D20626C616E64697420656C656D656E74756D206D61757269732C20766974;
        inPKT[126]      = 272'hC77E616520656C656D656E74756D20646F6C6F722068656E64726572697420766974;
        inPKT[127]      = 272'hC77F61652E204675736365206D6F6C65737469652C20656C697420757420616C6971;
        inPKT[128]      = 272'hC78075657420766F6C75747061742C206E657175652076656C697420707265746975;
        inPKT[129]      = 272'hC7816D2061756775652C206672696E67696C6C6120636F6E64696D656E74756D206A;
        inPKT[130]      = 272'hC7827573746F2073617069656E2061206A7573746F2E2050686173656C6C75732071;
        inPKT[131]      = 272'hC78375697320617563746F72206C6F72656D2C20696E20616C697175616D206E756E;
        inPKT[132]      = 272'hC784632E20557420656C656966656E6420616E7465206574206E697369206D6F6C65;
        inPKT[133]      = 272'hC7857374696520636F6E76616C6C69732069642065742073656D2E20536564206163;
        inPKT[134]      = 272'hC78620626962656E64756D20617263752E20467573636520766573746962756C756D;
        inPKT[135]      = 272'hC787206E756E6320656765742074656C6C7573206665726D656E74756D2C206E6563;
        inPKT[136]      = 272'hC7882072686F6E637573206D6173736120636F6D6D6F646F2E204D616563656E6173;
        inPKT[137]      = 272'hC789206964206E756E63206E6F6E20657820766573746962756C756D206F726E6172;
        inPKT[138]      = 272'hC78A65207574206E65632065726F732E20416C697175616D20656666696369747572;
        inPKT[139]      = 272'hC78B20636F6D6D6F646F206469616D206964206C6F626F727469732E205365642061;
        inPKT[140]      = 272'hC78C632074656D706F72206C65637475732E204E756E6320656C656D656E74756D20;
        inPKT[141]      = 272'hC78D7574206C65637475732061632074696E636964756E742E20557420696163756C;
        inPKT[142]      = 272'hC78E6973206E756C6C61207175697320657820656C656D656E74756D2C20616C6971;
        inPKT[143]      = 272'hC78F7565742073656D706572206D61676E6120656C656966656E642E0D0A0D0A4375;
        inPKT[144]      = 272'hC7907261626974757220746F72746F72206E69736C2C20756C747269636965732069;
        inPKT[145]      = 272'hC7916E206E657175652061632C20616363756D73616E20636F6E736571756174206D;
        inPKT[146]      = 272'hC792657475732E204D616563656E6173206D617373612073617069656E2C206D6174;
        inPKT[147]      = 272'hC79374697320696E2076656E656E617469732073697420616D65742C20617563746F;
        inPKT[148]      = 272'hC794722073697420616D657420656E696D2E204E756E63207669746165206D657475;
        inPKT[149]      = 272'hC7957320636F6D6D6F646F2C206D6174746973206D617373612073697420616D6574;
        inPKT[150]      = 272'hC7962C20766172697573206C6F72656D2E204E756E6320696E20656C697420656C69;
        inPKT[151]      = 272'hC797742E204E756E63206F726E61726520636F6E7365637465747572206D61676E61;
        inPKT[152]      = 272'hC7982C2073697420616D657420706F72747469746F7220617263752072686F6E6375;
        inPKT[153]      = 272'hC799732065752E2053757370656E6469737365207363656C6572697371756520756C;
        inPKT[154]      = 272'hC79A74726963696573206578206120616C697175616D2E2053757370656E64697373;
        inPKT[155]      = 272'hC79B652072757472756D20736F6C6C696369747564696E206E756E632C206E6F6E20;
        inPKT[156]      = 272'hC79C636F6E76616C6C697320747572706973206C616F726565742073697420616D65;
        inPKT[157]      = 272'hC79D742E2041656E65616E20612066696E69627573206D61757269732C2071756973;
        inPKT[158]      = 272'hC79E20637572737573206E756E632E20496E2066657567696174206475692076656C;
        inPKT[159]      = 272'hC79F2075726E612073656D7065722066617563696275732E204D617572697320756C;
        inPKT[160]      = 272'hC7A0747269636965732061742074757270697320656765742070656C6C656E746573;
        inPKT[161]      = 272'hC7A17175652E205072616573656E742073697420616D6574206C6967756C6120636F;
        inPKT[162]      = 272'hC7A26E76616C6C69732C20656C656D656E74756D206E756C6C6120756C6C616D636F;
        inPKT[163]      = 272'hC7A3727065722C20616C697175616D2075726E612E20457469616D207175616D2065;
        inPKT[164]      = 272'hC7A46C69742C20706F7375657265207574207175616D20656765742C2066696E6962;
        inPKT[165]      = 272'hC7A5757320736F6C6C696369747564696E206E756C6C612E20496E20737573636970;
        inPKT[166]      = 272'hC7A6697420656E696D2065742065726F732066696E696275732C207574207363656C;
        inPKT[167]      = 272'hC7A7657269737175652074656C6C757320666575676961742E204375726162697475;
        inPKT[168]      = 272'hC7A872206E6F6E206D617373612076617269757320646F6C6F722067726176696461;
        inPKT[169]      = 272'hC7A920656C656D656E74756D20717569732075742066656C69732E2050686173656C;
        inPKT[170]      = 272'hC7AA6C757320657569736D6F6420697073756D20656765742076656C6974206C6F62;
        inPKT[171]      = 272'hC7AB6F727469732C206567657420706F727461206D61757269732074656D7075732E;
        inPKT[172]      = 272'hC7AC2053656420696D7065726469657420766F6C75747061742074656C6C75732065;
        inPKT[173]      = 272'hC7AD752074696E636964756E742E0D0A0D0A55742076656C206D69206174206D6574;
        inPKT[174]      = 272'hC7AE7573206672696E67696C6C6120677261766964612E205072616573656E742065;
        inPKT[175]      = 272'hC7AF726F73206E6962682C2063757273757320656765737461732074696E63696475;
        inPKT[176]      = 272'hC7B06E7420736F64616C65732C207363656C65726973717565206E65632066656C69;
        inPKT[177]      = 272'hC7B1732E20496E746567657220696D70657264696574206D616C657375616461206E;
        inPKT[178]      = 272'hC7B269736C20616C69717565742076656E656E617469732E20496E74656765722073;
        inPKT[179]      = 272'hC7B3656420706F72747469746F7220697073756D2E20496E746567657220636F6D6D;
        inPKT[180]      = 272'hC7B46F646F206665756769617420746F72746F722C206575206C6F626F7274697320;
        inPKT[181]      = 272'hC7B5617567756520656C656D656E74756D2073697420616D65742E20446F6E656320;
        inPKT[182]      = 272'hC7B6766573746962756C756D206C6967756C612061756775652C2065742066696E69;
        inPKT[183]      = 272'hC7B7627573206172637520706F72746120696E2E204E756C6C612073656D2074656C;
        inPKT[184]      = 272'hC7B86C75732C20756C6C616D636F727065722061742063757273757320612C20706F;
        inPKT[185]      = 272'hC7B97274612073697420616D6574206D61676E612E204E756E632076697461652069;
        inPKT[186]      = 272'hC7BA6D706572646965742070757275732C206E656320736F6C6C696369747564696E;
        inPKT[187]      = 272'hC7BB2074656C6C75732E20416C697175616D206572617420766F6C75747061742E20;
        inPKT[188]      = 272'hC7BC536564206964206D61676E6120636F6D6D6F646F2C206C75637475732076656C;
        inPKT[189]      = 272'hC7BD697420717569732C20657569736D6F6420656E696D2E20496E7465676572206D;
        inPKT[190]      = 272'hC7BE617474697320736F64616C6573206665726D656E74756D2E2051756973717565;
        inPKT[191]      = 272'hC7BF20736564206672696E67696C6C61206C6F72656D2E2043726173207665686963;
        inPKT[192]      = 272'hC7C0756C612074656D7075732073617069656E20757420636F6E6775652E20447569;
        inPKT[193]      = 272'hC7C1732073617069656E20656E696D2C20706F727461206E6563206C656F2069642C;
        inPKT[194]      = 272'hC7C22065666669636974757220706F7375657265206C696265726F2E204E756C6C61;
        inPKT[195]      = 272'hC7C36D2061632074656D706F72206D657475732E205365642076656C207475727069;
        inPKT[196]      = 272'hC7C47320666575676961742C20696163756C697320617567756520717569732C2074;
        inPKT[197]      = 272'hC7C5696E636964756E74207475727069732E0D0A0D0A566976616D757320706F7375;
        inPKT[198]      = 272'hC7C665726520706F72747469746F722061756775652C207661726975732061636375;
        inPKT[199]      = 272'hC7C76D73616E20656C69742076756C70757461746520656765742E20517569737175;
        inPKT[200]      = 272'hC7C86520736564206D616C657375616461206E69736C2E20496E74657264756D2065;
        inPKT[201]      = 272'hC7C974206D616C6573756164612066616D657320616320616E746520697073756D20;
        inPKT[202]      = 272'hC7CA7072696D697320696E2066617563696275732E204E756E632074757270697320;
        inPKT[203]      = 272'hC7CB6469616D2C2073757363697069742061632065726F732076656C2C2074656D70;
        inPKT[204]      = 272'hC7CC75732076656E656E6174697320697073756D2E2044756973206C756374757320;
        inPKT[205]      = 272'hC7CD72686F6E637573206D617373612E204675736365207574206C6163696E696120;
        inPKT[206]      = 272'hC7CE7475727069732E20566976616D75732072757472756D2074656C6C7573206175;
        inPKT[207]      = 272'hC7CF6775652C206174206F726E617265206E69736C20666163696C69736973206574;
        inPKT[208]      = 272'hC7D02E204E756E6320736564206E6973692072697375732E20496E74656765722065;
        inPKT[209]      = 272'hC7D16C656D656E74756D206D6175726973207175616D2C207574207665686963756C;
        inPKT[210]      = 272'hC7D261206D617572697320636F6E6775652065752E0D0A0D0A467573636520612074;
        inPKT[211]      = 272'hC7D3656C6C75732073697420616D65742065726174206665726D656E74756D207363;
        inPKT[212]      = 272'hC7D4656C657269737175652E2043757261626974757220696E2076656C6974206174;
        inPKT[213]      = 272'hC7D520656E696D206C6163696E6961207665686963756C61206163206964206A7573;
        inPKT[214]      = 272'hC7D6746F2E2050726F696E206E6F6E20646F6C6F72206566666963697475722C2074;
        inPKT[215]      = 272'hC7D7696E636964756E74206F64696F2065752C20666175636962757320656E696D2E;
        inPKT[216]      = 272'hC7D82050656C6C656E7465737175652064617069627573206F726369206163206C6F;
        inPKT[217]      = 272'hC7D972656D20696163756C69732C2073697420616D657420626C616E646974206172;
        inPKT[218]      = 272'hC7DA6375207472697374697175652E2041656E65616E207472697374697175652074;
        inPKT[219]      = 272'hC7DB6F72746F72206E6563206A7573746F20616C697175616D2C20696E2070726574;
        inPKT[220]      = 272'hC7DC69756D2066656C6973206D6F6C65737469652E205365642065742074656D7075;
        inPKT[221]      = 272'hC7DD732061756775652E204E756C6C61206672696E67696C6C6120656C656966656E;
        inPKT[222]      = 272'hC7DE6420697073756D2076697665727261206375727375732E20416C697175616D20;
        inPKT[223]      = 272'hC7DF6D6178696D7573206665726D656E74756D206E69626820616320616363756D73;
        inPKT[224]      = 272'hC7E0616E2E204E756C6C6120666163696C6973692E20566573746962756C756D2066;
        inPKT[225]      = 272'hC7E16163696C69736973206C656F20656765737461732073656D206D617474697320;
        inPKT[226]      = 272'hC7E2636F6E6775652E204D6175726973207669746165206578206174207269737573;
        inPKT[227]      = 272'hC7E3206461706962757320656C656966656E642E20496E7465676572207574206572;
        inPKT[228]      = 272'hC7E46F7320636F6E6775652C20706F72747469746F7220616E7465206E6F6E2C2069;
        inPKT[229]      = 272'hC7E56E74657264756D20646F6C6F722E0D0A0D0A566573746962756C756D20656C65;
        inPKT[230]      = 272'hC7E66966656E64206D6175726973206575206E6973692064696374756D2067726176;
        inPKT[231]      = 272'hC7E76964612E2044756973206D6F6C6C6973206469616D2076656C20656E696D2074;
        inPKT[232]      = 272'hC7E8656D7075732C2076697461652064617069627573206D61737361207361676974;
        inPKT[233]      = 272'hC7E97469732E204E756C6C6120757420617563746F7220746F72746F722E204D6F72;
        inPKT[234]      = 272'hC7EA626920736564206C6F72656D2075726E612E204675736365206D61747469732C;
        inPKT[235]      = 272'hC7EB206D61676E6120616320636F6E64696D656E74756D20666575676961742C206D;
        inPKT[236]      = 272'hC7EC6173736120647569206D6178696D7573206E756C6C612C20657520616C697175;
        inPKT[237]      = 272'hC7ED6574206E65717565206D6175726973206120657261742E205175697371756520;
        inPKT[238]      = 272'hC7EE617563746F722065737420757420696E74657264756D20636F6E736563746574;
        inPKT[239]      = 272'hC7EF75722E20446F6E65632065676574206469676E697373696D20746F72746F722C;
        inPKT[240]      = 272'hC7F02068656E647265726974206D617474697320657261742E2050656C6C656E7465;
        inPKT[241]      = 272'hC7F173717565206861626974616E74206D6F72626920747269737469717565207365;
        inPKT[242]      = 272'hC7F26E6563747573206574206E65747573206574206D616C6573756164612066616D;
        inPKT[243]      = 272'hC7F365732061632074757270697320656765737461732E2051756973717565206F72;
        inPKT[244]      = 272'hC7F46E617265207661726975732074656D7075732E0D0A0D0A4D6F72626920727574;
        inPKT[245]      = 272'hC7F572756D20616E7465206E6962682C20612076697665727261206E756C6C612068;
        inPKT[246]      = 272'hC7F6656E64726572697420696E2E2050726F696E2073757363697069742065676573;
        inPKT[247]      = 272'hC7F774617320657261742C20757420617563746F72206F726369206D617474697320;
        inPKT[248]      = 272'hC7F8612E2050656C6C656E746573717565206C7563747573206672696E67696C6C61;
        inPKT[249]      = 272'hC7F920656C6974207574206C6163696E69612E205574206574206D61737361206E75;
        inPKT[250]      = 272'hC7FA6C6C612E20536564206174206672696E67696C6C61206C6F72656D2E2050726F;
        inPKT[251]      = 272'hC7FB696E206772617669646120616363756D73616E20726973757320736564206269;
        inPKT[252]      = 272'hC7FC62656E64756D2E204D616563656E6173206D616C657375616461206F64696F20;
        inPKT[253]      = 272'hC7FD75742076656C697420657569736D6F6420646170696275732E0D0A0D0A457469;
        inPKT[254]      = 272'hC7FE616D20636F6E677565206D617474697320696163756C69732E204D6175726973;
        inPKT[255]      = 272'hC7FF207669746165206566666963697475722073656D2E205365642070756C76696E;
        inPKT[256]      = 272'hC700617220646F6C6F72207574206D6920657569736D6F642068656E647265726974;
        inPKT[257]      = 272'hC7012E204E756C6C616D206174206772617669646120646F6C6F722E204D6F726269;
        inPKT[258]      = 272'hC702206C656F207475727069732C20636F6E677565206E656320616C697175616D20;
        inPKT[259]      = 272'hC70375742C20636F6D6D6F646F20696E206E756E632E204E756C6C61206174206661;
        inPKT[260]      = 272'hC704756369627573206C656F2C2065752066657567696174206C616375732E204675;
        inPKT[261]      = 272'hC705736365206E6F6E2065676573746173207475727069732E205175697371756520;
        inPKT[262]      = 272'hC706766974616520697073756D206D692E204E756E63206E6F6E206F726369207369;
        inPKT[263]      = 272'hC7077420616D6574206E6973692076617269757320706F72747469746F7220696E20;
        inPKT[264]      = 272'hC70876756C70757461746520746F72746F722E204E756E6320636F6E76616C6C6973;
        inPKT[265]      = 272'hC7092067726176696461206469616D206120756C747269636965732E205175697371;
        inPKT[266]      = 272'hC70A7565206575206A7573746F20636F6E64696D656E74756D2C2076617269757320;
        inPKT[267]      = 272'hC70B6469616D2076656C2C20766573746962756C756D206D617373612E0D0A0D0A50;
        inPKT[268]      = 272'hC70C656C6C656E7465737175652070656C6C656E7465737175652073617069656E20;
        inPKT[269]      = 272'hC70D6E657175652C20617563746F72206D616C65737561646120657261742068656E;
        inPKT[270]      = 272'hC70E647265726974206E65632E204E756C6C6120706C616365726174206469616D20;
        inPKT[271]      = 272'hC70F68656E647265726974206D6173736120626962656E64756D2C2061206D6F6C65;
        inPKT[272]      = 272'hC710737469652066656C69732068656E6472657269742E204D617572697320657569;
        inPKT[273]      = 272'hC711736D6F642076656E656E61746973206A7573746F2C20757420617563746F7220;
        inPKT[274]      = 272'hC712656C697420616C69717565742075742E20467573636520616C69717565742C20;
        inPKT[275]      = 272'hC7137175616D207574206469676E697373696D2068656E6472657269742C206D6175;
        inPKT[276]      = 272'hC71472697320747572706973206469676E697373696D20746F72746F722C20656765;
        inPKT[277]      = 272'hC715742070656C6C656E7465737175652076656C6974206F726369206E6563207175;
        inPKT[278]      = 272'hC716616D2E204E756E6320656765737461732070656C6C656E746573717565207269;
        inPKT[279]      = 272'hC7177375732E204375726162697475722073757363697069742074656D707573206C;
        inPKT[280]      = 272'hC718616375732C2065676574207072657469756D20656C69742074696E636964756E;
        inPKT[281]      = 272'hC71974206E6F6E2E20437261732075726E61206C6F72656D2C20706C616365726174;
        inPKT[282]      = 272'hC71A20766F6C757470617420696D706572646965742073697420616D65742C206567;
        inPKT[283]      = 272'hC71B65737461732076656C206F7263692E0D0A0D0A50656C6C656E74657371756520;
        inPKT[284]      = 272'hC71C736F64616C6573206665726D656E74756D206E69736C2C206174206672696E67;
        inPKT[285]      = 272'hC71D696C6C61206475692073656D706572206665726D656E74756D2E204E756C6C61;
        inPKT[286]      = 272'hC71E6D20706C6163657261742076656C206D692068656E64726572697420656C656D;
        inPKT[287]      = 272'hC71F656E74756D2E20457469616D206E6F6E20697073756D2065782E204E616D2061;
        inPKT[288]      = 272'hC72063207363656C65726973717565206E6962682C2076656C20666163696C697369;
        inPKT[289]      = 272'hC72173206D692E20446F6E65632065676573746173206C616F726565742065726F73;
        inPKT[290]      = 272'hC7222C206567657420766F6C7574706174206D657475732E205072616573656E7420;
        inPKT[291]      = 272'hC723616363756D73616E20626962656E64756D206E69736C206E65632076656E656E;
        inPKT[292]      = 272'hC724617469732E205365642072757472756D206D6920612073757363697069742070;
        inPKT[293]      = 272'hC725686172657472612E205365642073697420616D657420696E74657264756D2074;
        inPKT[294]      = 272'hC72675727069732E20416C697175616D206575206E69626820746F72746F722E2044;
        inPKT[295]      = 272'hC7276F6E65632066617563696275732064617069627573206E6973692C2073656420;
        inPKT[296]      = 272'hC7286C616F72656574206F726369207363656C6572697371756520696E2E0D0A0D0A;
        inPKT[297]      = 272'hC7294D617572697320696E2066656C6973206665726D656E74756D2C20636F6E7661;
        inPKT[298]      = 272'hC72A6C6C69732061756775652076656C2C20706F7375657265206D692E2050656C6C;
        inPKT[299]      = 272'hC72B656E746573717565207363656C657269737175652072686F6E637573206A7573;
        inPKT[300]      = 272'hC72C746F2C2065752070756C76696E617220656E696D2070756C76696E6172207665;
        inPKT[301]      = 272'hC72D6C2E204D616563656E6173207068617265747261206C696265726F206D61676E;
        inPKT[302]      = 272'hC72E612C20616320736F6C6C696369747564696E206C656F206D6F6C6C6973206E6F;
        inPKT[303]      = 272'hC72F6E2E204E756C6C6120656C656D656E74756D206F726E61726520656765737461;
        inPKT[304]      = 272'hC730732E20436C61737320617074656E742074616369746920736F63696F73717520;
        inPKT[305]      = 272'hC7316164206C69746F726120746F727175656E742070657220636F6E75626961206E;
        inPKT[306]      = 272'hC7326F737472612C2070657220696E636570746F732068696D656E61656F732E2050;
        inPKT[307]      = 272'hC73372616573656E74206175677565206D61757269732C2072686F6E637573207175;
        inPKT[308]      = 272'hC734697320657374206E6F6E2C206D6F6C6C697320636F6E76616C6C69732066656C;
        inPKT[309]      = 272'hC73569732E2053757370656E646973736520666163696C697369732C206F72636920;
        inPKT[310]      = 272'hC7367669746165206C6163696E69612074656D706F722C206C656374757320736170;
        inPKT[311]      = 272'hC73769656E206D61747469732072697375732C206E6F6E2073616769747469732065;
        inPKT[312]      = 272'hC7386C6974206E657175652071756973206A7573746F2E20446F6E6563206D616C65;
        inPKT[313]      = 272'hC7397375616461206C6163696E6961206475692E2050686173656C6C75732068656E;
        inPKT[314]      = 272'hC73A647265726974206D6175726973206D61757269732C20736564206672696E6769;
        inPKT[315]      = 272'hC73B6C6C61206C696265726F206672696E67696C6C6120696E2E2053656420617420;
        inPKT[316]      = 272'hC73C6C6967756C6120696E206A7573746F2066696E696275732076756C7075746174;
        inPKT[317]      = 272'hC73D652E204E756E6320637572737573206E657175652073697420616D6574206172;
        inPKT[318]      = 272'hC73E63752074696E636964756E742C2076697461652070686172657472612073656D;
        inPKT[319]      = 272'hC73F20706F72747469746F722E20416C697175616D206D61747469732C206A757374;
        inPKT[320]      = 272'hC7406F206E6F6E20657569736D6F6420636F6E76616C6C69732C206E756E63206D69;
        inPKT[321]      = 272'hC74120636F6E736571756174206573742C206E656320736F6C6C696369747564696E;
        inPKT[322]      = 272'hC742206C65637475732073617069656E2076656C206F64696F2E20496E2074656D70;
        inPKT[323]      = 272'hC7436F72206572617420646F6C6F722C20736564207665686963756C612075726E61;
        inPKT[324]      = 272'hC74420636F6E736571756174207365642E0D0A0D0A4E616D2072686F6E6375732069;
        inPKT[325]      = 272'hC74564206D6175726973206E6563206469676E697373696D2E20496E20696D706572;
        inPKT[326]      = 272'hC7466469657420756C7472696365732065726174206E656320736F6C6C6963697475;
        inPKT[327]      = 272'hC74764696E2E20496E74656765722073656420636F6E64696D656E74756D2065726F;
        inPKT[328]      = 272'hC748732E20446F6E65632065676574206E756E63206964206D617572697320747269;
        inPKT[329]      = 272'hC74973746971756520706F72747469746F72206C616F72656574207669746165206D;
        inPKT[330]      = 272'hC74A657475732E204E756C6C6120666163696C6973692E204E756C6C616D20657520;
        inPKT[331]      = 272'hC74B6C616375732061206469616D207472697374697175652065676573746173206E;
        inPKT[332]      = 272'hC74C6F6E20696163756C6973206D657475732E20416C697175616D20696E2074656D;
        inPKT[333]      = 272'hC74D706F7220657261742C20696420636F6E677565206D617373612E20566976616D;
        inPKT[334]      = 272'hC74E75732076656C20746F72746F72207669746165206E69626820636F6D6D6F646F;
        inPKT[335]      = 272'hC74F206C6F626F727469732071756973206120697073756D2E2050726F696E20766F;
        inPKT[336]      = 272'hC7506C7574706174207175616D206E6F6E2066656C69732074656D7075732C206964;
        inPKT[337]      = 272'hC75120706F737565726520646F6C6F722074656D706F722E205072616573656E7420;
        inPKT[338]      = 272'hC75276697461652074696E636964756E742073617069656E2E204D616563656E6173;
        inPKT[339]      = 272'hC75320666163696C69736973206D617474697320616E746520717569732076617269;
        inPKT[340]      = 272'hC75475732E20446F6E65632070656C6C656E7465737175652065726F732066657567;
        inPKT[341]      = 272'hC7556961742074696E636964756E7420636F6E64696D656E74756D2E2050726F696E;
        inPKT[342]      = 272'hC75620666175636962757320766F6C7574706174206D692073656420736167697474;
        inPKT[343]      = 272'hC75769732E0D0A0D0A44756973206772617669646120656C656D656E74756D20696E;
        inPKT[344]      = 272'hC75874657264756D2E2050726F696E2073697420616D6574207175616D206C696775;
        inPKT[345]      = 272'hC7596C612E2050686173656C6C757320636F6D6D6F646F2C2075726E6120696E2063;
        inPKT[346]      = 272'hC75A6F6E67756520766F6C75747061742C206C6967756C6120657820706861726574;
        inPKT[347]      = 272'hC75B7261206C6967756C612C20696E2064696374756D206D61676E61206F72636920;
        inPKT[348]      = 272'hC75C6E6563206D61757269732E204E756E6320617563746F7220636F6E7365637465;
        inPKT[349]      = 272'hC75D74757220766F6C75747061742E204D6F7262692074696E636964756E74206E69;
        inPKT[350]      = 272'hC75E626820757420656E696D2065666669636974757220677261766964612E204375;
        inPKT[351]      = 272'hC75F72616269747572207669746165207175616D2065726F732E2044756973206672;
        inPKT[352]      = 272'hC760696E67696C6C6120616320746F72746F7220696E2074696E636964756E742E20;
        inPKT[353]      = 272'hC7614E756E632076656C206D61757269732072697375732E20446F6E656320656C65;
        inPKT[354]      = 272'hC7626966656E64206C6967756C61207361676974746973206E6973692066696E6962;
        inPKT[355]      = 272'hC76375732C2061207363656C65726973717565206C696265726F2070656C6C656E74;
        inPKT[356]      = 272'hC76465737175652E20566573746962756C756D20747269737469717565206D617373;
        inPKT[357]      = 272'hC76561206E6962682C20617420766573746962756C756D206D61676E612066696E69;
        inPKT[358]      = 272'hC7666275732065752E0D0A0D0A43757261626974757220696D706572646965742070;
        inPKT[359]      = 272'hC767757275732065676574206E756E6320756C7472696365732C2076697461652076;
        inPKT[360]      = 272'hC768656E656E61746973206D6173736120636F6D6D6F646F2E2050656C6C656E7465;
        inPKT[361]      = 272'hC76973717565206861626974616E74206D6F72626920747269737469717565207365;
        inPKT[362]      = 272'hC76A6E6563747573206574206E65747573206574206D616C6573756164612066616D;
        inPKT[363]      = 272'hC76B65732061632074757270697320656765737461732E20496E206665726D656E74;
        inPKT[364]      = 272'hC76C756D2061742075726E61206E6F6E20636F6E76616C6C69732E20446F6E656320;
        inPKT[365]      = 272'hC76D6163206175677565206A7573746F2E20496E20617420656C6974206574206172;
        inPKT[366]      = 272'hC76E6375206D6178696D7573206C75637475732E20467573636520657569736D6F64;
        inPKT[367]      = 272'hC76F206E756E63206E65632076656E656E6174697320617563746F722E204C6F7265;
        inPKT[368]      = 272'hC7706D20697073756D20646F6C6F722073697420616D65742C20636F6E7365637465;
        inPKT[369]      = 272'hC7717475722061646970697363696E6720656C69742E20446F6E6563206469637475;
        inPKT[370]      = 272'hC7726D2074656D706F722072757472756D2E2053656420656C656966656E64206469;
        inPKT[371]      = 272'hC773616D206964206D6173736120696D706572646965742C206163206F726E617265;
        inPKT[372]      = 272'hC774206C696265726F20656C656966656E642E204D616563656E6173206F726E6172;
        inPKT[373]      = 272'hC77565206D65747573206E756C6C612C2073697420616D6574206665726D656E7475;
        inPKT[374]      = 272'hC7766D20656C697420616C697175616D2069642E20446F6E656320756C7472696365;
        inPKT[375]      = 272'hC7777320746F72746F7220617420616E74652068656E6472657269742C2065752073;
        inPKT[376]      = 272'hC77861676974746973206A7573746F20756C7472696365732E0D0A0D0A5072616573;
        inPKT[377]      = 272'hC779656E74206C7563747573207072657469756D206E657175652C2073697420616D;
        inPKT[378]      = 272'hC77A65742070656C6C656E746573717565206D617572697320656C656D656E74756D;
        inPKT[379]      = 272'hC77B206E6F6E2E20557420626C616E646974207068617265747261206F64696F206E;
        inPKT[380]      = 272'hC77C6F6E20657569736D6F642E2051756973717565207669746165206C656F20616C;
        inPKT[381]      = 272'hC77D697175616D2C20736F64616C65732074656C6C75732069642C20696163756C69;
        inPKT[382]      = 272'hC77E73206D61757269732E204E616D2065666669636974757220696E207075727573;
        inPKT[383]      = 272'hC77F2073656420616363756D73616E2E204D616563656E61732073697420616D6574;
        inPKT[384]      = 272'hC780206375727375732066656C69732E20517569737175652066617563696275732C;
        inPKT[385]      = 272'hC7812064756920657420617563746F72206C75637475732C20616E74652065726174;
        inPKT[386]      = 272'hC78220706F73756572652065726F732C20757420636F6E76616C6C6973206D657475;
        inPKT[387]      = 272'hC78373206C6563747573207669746165206C656F2E2053757370656E646973736520;
        inPKT[388]      = 272'hC784706F74656E74692E204372617320657420646F6C6F72206E6F6E2075726E6120;
        inPKT[389]      = 272'hC7857363656C65726973717565207472697374697175652E20437261732072757472;
        inPKT[390]      = 272'hC786756D206E65632076656C69742061632073616769747469732E20446F6E656320;
        inPKT[391]      = 272'hC787656C656966656E642C206C61637573207365642067726176696461206D616C65;
        inPKT[392]      = 272'hC78873756164612C20657820616E746520706C616365726174206C65637475732C20;
        inPKT[393]      = 272'hC7896567657420636F6E677565206D61737361206D65747573206964206C61637573;
        inPKT[394]      = 272'hC78A2E2053757370656E64697373652069642072757472756D206C65637475732E20;
        inPKT[395]      = 272'hC78B4675736365206D6178696D757320736564206C6967756C612073656420766976;
        inPKT[396]      = 272'hC78C657272612E204E616D206C7563747573206469616D20616E74652C2076697461;
        inPKT[397]      = 272'hC78D65206F726E617265206E657175652076617269757320656765742E0D0A0D0A50;
        inPKT[398]      = 272'hC78E656C6C656E74657371756520617420656C6974206E6962682E20566573746962;
        inPKT[399]      = 272'hC78F756C756D20616E746520697073756D207072696D697320696E20666175636962;
        inPKT[400]      = 272'hC7907573206F726369206C756374757320657420756C74726963657320706F737565;
        inPKT[401]      = 272'hC791726520637562696C69612043757261653B204375726162697475722066617563;
        inPKT[402]      = 272'hC79269627573206469616D206C656F2C206E656320657569736D6F642073656D2065;
        inPKT[403]      = 272'hC79366666963697475722075742E205574207665686963756C612061756775652061;
        inPKT[404]      = 272'hC79463206C696265726F20696163756C69732C206E656320656C656966656E642065;
        inPKT[405]      = 272'hC7957820706F7274612E204D6F7262692068656E6472657269742067726176696461;
        inPKT[406]      = 272'hC7962074696E636964756E742E205072616573656E7420646F6C6F72206C61637573;
        inPKT[407]      = 272'hC7972C2074656D707573206575206672696E67696C6C612073697420616D65742C20;
        inPKT[408]      = 272'hC798656C656966656E6420696E206E756C6C612E204E756C6C61206D6F6C6C697320;
        inPKT[409]      = 272'hC79965676574206D61676E61206E65632068656E6472657269742E20416C69717561;
        inPKT[410]      = 272'hC79A6D20636F6E76616C6C69732073656D2076697461652073617069656E20646963;
        inPKT[411]      = 272'hC79B74756D2C20757420766573746962756C756D206C6F72656D206672696E67696C;
        inPKT[412]      = 272'hC79C6C612E20446F6E65632074656C6C7573206C696265726F2C2066657567696174;
        inPKT[413]      = 272'hC79D2075742066696E69627573206E65632C20616C697175616D2073697420616D65;
        inPKT[414]      = 272'hC79E74206F7263692E204E756E63207375736369706974206E69736C206574206F72;
        inPKT[415]      = 272'hC79F6E61726520766573746962756C756D2E204E756C6C616D206C6F626F72746973;
        inPKT[416]      = 272'hC7A02073617069656E206A7573746F2C2073697420616D6574206469676E69737369;
        inPKT[417]      = 272'hC7A16D206E756C6C6120636F6E64696D656E74756D20696E2E20536564206D6F6C65;
        inPKT[418]      = 272'hC7A27374696520766F6C7574706174206E697369206174206665726D656E74756D2E;
        inPKT[419]      = 272'hC7A3204E756C6C61206D6F6C6573746965206E697369207365642074757270697320;
        inPKT[420]      = 272'hC7A46D6F6C65737469652C206E6F6E20696163756C6973206E756E63206661756369;
        inPKT[421]      = 272'hC7A56275732E2041656E65616E20696E74657264756D20706861726574726120636F;
        inPKT[422]      = 272'hC7A66E73656374657475722E20457469616D206578206F7263692C20696163756C69;
        inPKT[423]      = 272'hC7A773206E6F6E20657569736D6F642069642C20756C6C616D636F72706572207363;
        inPKT[424]      = 272'hC7A8656C65726973717565206F64696F2E0D0A0D0A4E616D20756C74726963657320;
        inPKT[425]      = 272'hC7A9656C656966656E64206469616D2C206567657420736F64616C65732073656D20;
        inPKT[426]      = 272'hC7AA6D61747469732061632E2055742076656E656E61746973206E69626820657520;
        inPKT[427]      = 272'hC7AB6C65637475732074696E636964756E742064696374756D2E20566976616D7573;
        inPKT[428]      = 272'hC7AC206375727375732061756775652071756973206C6F626F727469732065756973;
        inPKT[429]      = 272'hC7AD6D6F642E204E756E6320616C697175616D206469616D20617420616E74652066;
        inPKT[430]      = 272'hC7AE6163696C69736973206D6178696D75732E20457469616D20736564206C6F7265;
        inPKT[431]      = 272'hC7AF6D206D61747469732C20636F6E76616C6C69732075726E612076697461652C20;
        inPKT[432]      = 272'hC7B074656D7075732073656D2E20566976616D7573206567657374617320766F6C75;
        inPKT[433]      = 272'hC7B1747061742065726F7320657520756C7472696365732E20566573746962756C75;
        inPKT[434]      = 272'hC7B26D20756C6C616D636F727065722065726174206E756E632C206E6F6E2068656E;
        inPKT[435]      = 272'hC7B3647265726974206F64696F2070656C6C656E7465737175652069642E20467573;
        inPKT[436]      = 272'hC7B463652075726E6120697073756D2C206C6163696E696120696E20737573636970;
        inPKT[437]      = 272'hC7B569742076656C2C2073656D70657220696E206F64696F2E2050656C6C656E7465;
        inPKT[438]      = 272'hC7B673717565206964206E696268206E6973692E20416C697175616D20706F727461;
        inPKT[439]      = 272'hC7B7206E69736C20657420657820696163756C6973207472697374697175652E2045;
        inPKT[440]      = 272'hC7B87469616D206D61737361206F7263692C206567657374617320736564206C6F72;
        inPKT[441]      = 272'hC7B9656D20717569732C206469676E697373696D2073656D70657220616E74652E20;
        inPKT[442]      = 272'hC7BA53757370656E64697373652074696E636964756E74206E6973692065782C2073;
        inPKT[443]      = 272'hC7BB656420766F6C757470617420657374207661726975732076697461652E0D0A0D;
        inPKT[444]      = 272'hC7BC0A5365642073656D706572206C6163696E696120646F6C6F722E204E616D2075;
        inPKT[445]      = 272'hC7BD742076656C697420696E206C6163757320636F6E736563746574757220636F6E;
        inPKT[446]      = 272'hC7BE76616C6C69732070656C6C656E746573717565207365642073656D2E20537573;
        inPKT[447]      = 272'hC7BF70656E646973736520636F6E64696D656E74756D20612065726F732069642075;
        inPKT[448]      = 272'hC7C06C6C616D636F727065722E204D6F726269206C75637475732075726E61207369;
        inPKT[449]      = 272'hC7C17420616D657420657569736D6F6420696163756C69732E2050656C6C656E7465;
        inPKT[450]      = 272'hC7C27371756520666163696C69736973206D617572697320657520656C656D656E74;
        inPKT[451]      = 272'hC7C3756D207661726975732E204F72636920766172697573206E61746F7175652070;
        inPKT[452]      = 272'hC7C4656E617469627573206574206D61676E6973206469732070617274757269656E;
        inPKT[453]      = 272'hC7C574206D6F6E7465732C206E61736365747572207269646963756C7573206D7573;
        inPKT[454]      = 272'hC7C62E20446F6E6563206469676E697373696D206120697073756D20756C74726963;
        inPKT[455]      = 272'hC7C76965732076656E656E617469732E20566976616D7573206E756E632076656C69;
        inPKT[456]      = 272'hC7C8742C207665686963756C61207669746165206D617373612075742C20636F6E76;
        inPKT[457]      = 272'hC7C9616C6C697320636F6E736563746574757220746F72746F722E20517569737175;
        inPKT[458]      = 272'hC7CA6520616C697175616D2C206E69736C20636F6E67756520626C616E6469742075;
        inPKT[459]      = 272'hC7CB6C747269636965732C2075726E6120747572706973206D6174746973206D6167;
        inPKT[460]      = 272'hC7CC6E612C206E6F6E206665726D656E74756D206475692076656C69742065752071;
        inPKT[461]      = 272'hC7CD75616D2E0D0A0D0A496E2070686172657472612076656C697420646F6C6F722C;
        inPKT[462]      = 272'hC7CE20766974616520637572737573206F7263692066696E696275732074696E6369;
        inPKT[463]      = 272'hC7CF64756E742E20566976616D757320696420746F72746F722072686F6E6375732C;
        inPKT[464]      = 272'hC7D0207361676974746973206469616D20656765742C207072657469756D206D6175;
        inPKT[465]      = 272'hC7D17269732E2050686173656C6C757320656C656D656E74756D20656E696D206665;
        inPKT[466]      = 272'hC7D26C69732E204D6175726973206575206E65717565206567657420707572757320;
        inPKT[467]      = 272'hC7D368656E64726572697420677261766964612E20416C697175616D206C69626572;
        inPKT[468]      = 272'hC7D46F206E6962682C20636F6E76616C6C69732061206E69736C2065742C2068656E;
        inPKT[469]      = 272'hC7D564726572697420766573746962756C756D2066656C69732E20446F6E65632065;
        inPKT[470]      = 272'hC7D67569736D6F64206665726D656E74756D2074757270697320657520617563746F;
        inPKT[471]      = 272'hC7D7722E2041656E65616E20626962656E64756D2074757270697320696E206F6469;
        inPKT[472]      = 272'hC7D86F20636F6E76616C6C69732C20766974616520766172697573206578206C616F;
        inPKT[473]      = 272'hC7D9726565742E2046757363652076656C206D6920766974616520646F6C6F722066;
        inPKT[474]      = 272'hC7DA6575676961742076756C707574617465206E6563207574206E756E632E204372;
        inPKT[475]      = 272'hC7DB617320646170696275732C20616E7465206964207665686963756C6120616C69;
        inPKT[476]      = 272'hC7DC7175616D2C20656C69742065726F73207361676974746973206D692C206E6F6E;
        inPKT[477]      = 272'hC7DD20656C656966656E64206578206E756C6C6120656765742076656C69742E2053;
        inPKT[478]      = 272'hC7DE757370656E6469737365206964206469616D206475692E2053757370656E6469;
        inPKT[479]      = 272'hC7DF737365207072657469756D206A7573746F20736564206E69626820706F727474;
        inPKT[480]      = 272'hC7E069746F722C2076656C20696E74657264756D206D6175726973206D6178696D75;
        inPKT[481]      = 272'hC7E1732E20557420616C697175616D206C616375732070757275732C207369742061;
        inPKT[482]      = 272'hC7E26D657420696D70657264696574206E69626820666575676961742069642E2049;
        inPKT[483]      = 272'hC7E36E7465676572206C6F72656D206D61757269732C207072657469756D206E6F6E;
        inPKT[484]      = 272'hC7E4206E6973692065742C20646170696275732066696E69627573206F7263692E0D;
        inPKT[485]      = 272'hC7E50A0D0A566573746962756C756D20696163756C69732C206D61676E6120617420;
        inPKT[486]      = 272'hC7E66D6174746973206D6178696D75732C2061726375206572617420646170696275;
        inPKT[487]      = 272'hC7E773206E756E632C206120766172697573206D657475732066656C697320736564;
        inPKT[488]      = 272'hC7E8206F7263692E204E756C6C616D206D69206E6962682C20656C656966656E6420;
        inPKT[489]      = 272'hC7E96E656320756C747269636573206E65632C20636F6E7365637465747572206163;
        inPKT[490]      = 272'hC7EA20656E696D2E20536564206C75637475732073656D20717569732074656D706F;
        inPKT[491]      = 272'hC7EB7220636F6E6775652E2053757370656E646973736520706F74656E74692E2045;
        inPKT[492]      = 272'hC7EC7469616D2065676574206C696265726F2076656C69742E204475697320766573;
        inPKT[493]      = 272'hC7ED746962756C756D20636F6E73657175617420706F7274612E204D617572697320;
        inPKT[494]      = 272'hC7EE706F72747469746F722074757270697320696E206D6173736120616C69717561;
        inPKT[495]      = 272'hC7EF6D20636F6E6775652E204E756C6C6120636F6E73656374657475722075726E61;
        inPKT[496]      = 272'hC7F0206D657475732C20696420696163756C6973206E756E6320756C747269636965;
        inPKT[497]      = 272'hC7F17320656765742E20437572616269747572206D6175726973206E657175652C20;
        inPKT[498]      = 272'hC7F2626962656E64756D207365642065726F732061742C206D6178696D757320756C;
        inPKT[499]      = 272'hC7F3747269636573207475727069732E0D0A496E74657264756D206574206D616C65;
        inPKT[500]      = 272'hC7F473756164612066616D657320616320616E746520697073756D207072696D6973;
        inPKT[501]      = 272'hC7F520696E2066617563696275732E2050656C6C656E74657371756520736F6C6C69;
        inPKT[502]      = 272'hC7F66369747564696E20626C616E646974206665726D656E74756D2E2050656C6C65;
        inPKT[503]      = 272'hC7F76E746573717565206E6F6E206C6967756C6120657520657261742076656E656E;
        inPKT[504]      = 272'hC7F86174697320657569736D6F642E2050656C6C656E74657371756520736F64616C;
        inPKT[505]      = 272'hC7F9657320766573746962756C756D20636F6E76616C6C69732E2050726F696E206D;
        inPKT[506]      = 272'hC7FA6F6C6573746965207072657469756D2065726F732076656C2065676573746173;
        inPKT[507]      = 272'hC7FB2E204D6F72626920736F6C6C696369747564696E207075727573206163206665;
        inPKT[508]      = 272'hC7FC726D656E74756D206D61747469732E204E756E632076656C2074696E63696475;
        inPKT[509]      = 272'hC7FD6E74206C696265726F2E204E756C6C6120616C697175657420697073756D206E;
        inPKT[510]      = 272'hC7FE6563207175616D20696D7065726469657420696E74657264756D2E2050726165;
        inPKT[511]      = 272'hC7FF73656E74206C6967756C612066656C69732C20696163756C697320617420616C;
        inPKT[512]      = 272'hC70069717565742061742C207361676974746973207175697320656C69742E0D0A51;
        inPKT[513]      = 272'hC7017569737175652076656C20696D70657264696574206E6962682E205068617365;
        inPKT[514]      = 272'hC7026C6C75732072757472756D206469676E697373696D207269737573206E6F6E20;
        inPKT[515]      = 272'hC70374696E636964756E742E20566573746962756C756D206E756E6320697073756D;
        inPKT[516]      = 272'hC7042C2076656E656E61746973206567657420706F72746120696E2C20636F6E7365;
        inPKT[517]      = 272'hC70563746574757220657520657261742E20446F6E6563207665686963756C612061;
        inPKT[518]      = 272'hC7066E74652076656C2072686F6E6375732066617563696275732E2050656C6C656E;
        inPKT[519]      = 272'hC707746573717565206A7573746F20746F72746F722C20766F6C757470617420696E;
        inPKT[520]      = 272'hC708206D61757269732061742C207661726975732070686172657472612072697375;
        inPKT[521]      = 272'hC709732E2051756973717565207574206469616D2073757363697069742C20736F6C;
        inPKT[522]      = 272'hC70A6C696369747564696E2073617069656E2065742C20696E74657264756D206C61;
        inPKT[523]      = 272'hC70B6375732E204D6F7262692072697375732073656D2C2070656C6C656E74657371;
        inPKT[524]      = 272'hC70C75652065742074757270697320696E2C20626C616E64697420736F6C6C696369;
        inPKT[525]      = 272'hC70D747564696E2073656D2E2053656420656666696369747572206C696265726F20;
        inPKT[526]      = 272'hC70E71756973207072657469756D207072657469756D2E204E756C6C616D20617563;
        inPKT[527]      = 272'hC70F746F72207361676974746973206C6F72656D2C20616320756C74726963657320;
        inPKT[528]      = 272'hC71061726375206D6178696D757320656765742E0D0A566573746962756C756D2076;
        inPKT[529]      = 272'hC7116F6C7574706174206C6967756C6120617563746F722073656D20766976657272;
        inPKT[530]      = 272'hC712612C20756C6C616D636F7270657220657569736D6F64206E6571756520706F72;
        inPKT[531]      = 272'hC713747469746F722E2053757370656E64697373652076697665727261207363656C;
        inPKT[532]      = 272'hC71465726973717565206F64696F2072686F6E63757320766F6C75747061742E2041;
        inPKT[533]      = 272'hC7156C697175616D206572617420766F6C75747061742E2053757370656E64697373;
        inPKT[534]      = 272'hC7166520706F74656E74692E20496E206861632068616269746173736520706C6174;
        inPKT[535]      = 272'hC71765612064696374756D73742E2050726F696E207574206E756C6C612075742064;
        inPKT[536]      = 272'hC7187569207363656C657269737175652064696374756D2E20517569737175652073;
        inPKT[537]      = 272'hC71975736369706974206E69626820706F7375657265207175616D2076756C707574;
        inPKT[538]      = 272'hC71A6174652C206575206C6163696E696120616E746520677261766964612E204375;
        inPKT[539]      = 272'hC71B72616269747572206D61737361206C6F72656D2C206F726E617265206575206D;
        inPKT[540]      = 272'hC71C6F6C6C69732061742C207068617265747261206E6563206D617373612E204E75;
        inPKT[541]      = 272'hC71D6C6C612066696E6962757320656C656966656E64206F7263692073697420616D;
        inPKT[542]      = 272'hC71E657420636F6E73656374657475722E205365642074656D707573207669746165;
        inPKT[543]      = 272'hC71F2061726375206E6563206665726D656E74756D2E2041656E65616E2070656C6C;
        inPKT[544]      = 272'hC720656E74657371756520766974616520646F6C6F7220696E20616363756D73616E;
        inPKT[545]      = 272'hC7212E2043726173206469676E697373696D2076756C707574617465206D6F6C6C69;
        inPKT[546]      = 272'hC722732E204D617572697320706F7274612076656E656E617469732072697375732C;
        inPKT[547]      = 272'hC7232065752074726973746971756520646F6C6F722072757472756D20696E2E2046;
        inPKT[548]      = 272'hC7247573636520636F6E64696D656E74756D206F7263692066656C69732C20736974;
        inPKT[549]      = 272'hC72520616D657420636F6E76616C6C6973206C696265726F2074696E636964756E74;
        inPKT[550]      = 272'hC7262061632E0D0A566573746962756C756D20696D7065726469657420656C697420;
        inPKT[551]      = 272'hC72774656D706F72207175616D20677261766964612C207574206D616C6573756164;
        inPKT[552]      = 272'hC728612074656C6C757320696D706572646965742E2050686173656C6C7573206F64;
        inPKT[553]      = 272'hC729696F2073656D2C206D61747469732073656420756C7472696365732061742C20;
        inPKT[554]      = 272'hC72A766976657272612076656C206475692E204E756E632075726E61206D65747573;
        inPKT[555]      = 272'hC72B2C206C7563747573206163206D6178696D757320696E2C20636F6E7365637465;
        inPKT[556]      = 272'hC72C747572206E6F6E206E6973692E204E756C6C612073697420616D657420626962;
        inPKT[557]      = 272'hC72D656E64756D2076656C69742E20446F6E6563207175697320656E696D206E6F6E;
        inPKT[558]      = 272'hC72E20726973757320626C616E64697420666163696C697369732071756973206E65;
        inPKT[559]      = 272'hC72F632072697375732E204375726162697475722065752065737420766974616520;
        inPKT[560]      = 272'hC7306C656374757320626C616E64697420616C69717565742E20566573746962756C;
        inPKT[561]      = 272'hC731756D20616E746520697073756D207072696D697320696E206661756369627573;
        inPKT[562]      = 272'hC732206F726369206C756374757320657420756C74726963657320706F7375657265;
        inPKT[563]      = 272'hC73320637562696C69612043757261653B20566573746962756C756D206163206469;
        inPKT[564]      = 272'hC734676E697373696D206E756E632E205175697371756520696E2073616769747469;
        inPKT[565]      = 272'hC735732074656C6C75732C2073697420616D6574206665726D656E74756D206E6962;
        inPKT[566]      = 272'hC736682E0D0A496E206469676E697373696D20726973757320766974616520707572;
        inPKT[567]      = 272'hC737757320766573746962756C756D2C20617420656C656D656E74756D206E756C6C;
        inPKT[568]      = 272'hC7386120706F73756572652E20536564206D6174746973206E756E63206E6962682E;
        inPKT[569]      = 272'hC7392053757370656E64697373652070656C6C656E74657371756520706C61636572;
        inPKT[570]      = 272'hC73A6174207363656C657269737175652E2041656E65616E2066657567696174206D;
        inPKT[571]      = 272'hC73B617572697320696420636F6E677565206C6163696E69612E20457469616D2073;
        inPKT[572]      = 272'hC73C75736369706974206C6967756C612074656C6C75732C206120636F6E67756520;
        inPKT[573]      = 272'hC73D6C656374757320616C697175616D207665686963756C612E2053757370656E64;
        inPKT[574]      = 272'hC73E69737365206567657420616E74652076656C20656E696D206D616C6573756164;
        inPKT[575]      = 272'hC73F6120766976657272612E2050726F696E2074696E636964756E74206172637520;
        inPKT[576]      = 272'hC740656765742076756C70757461746520616363756D73616E2E20496E2076697461;
        inPKT[577]      = 272'hC74165206469616D206E6962682E204D6F726269206D6178696D75732066656C6973;
        inPKT[578]      = 272'hC74220696420636F6E736563746574757220616C697175616D2E204E756C6C612066;
        inPKT[579]      = 272'hC7436163696C6973692E0D0A566573746962756C756D20766573746962756C756D20;
        inPKT[580]      = 272'hC74465666669636974757220746F72746F722073697420616D657420666163696C69;
        inPKT[581]      = 272'hC7457369732E204D616563656E6173206E6F6E2074656C6C7573206F7263692E2050;
        inPKT[582]      = 272'hC746686173656C6C7573206E6F6E206C7563747573206A7573746F2C206174207375;
        inPKT[583]      = 272'hC7477363697069742074656C6C75732E2046757363652068656E647265726974206E;
        inPKT[584]      = 272'hC7486563206E6962682076656C206375727375732E2053757370656E646973736520;
        inPKT[585]      = 272'hC749706F74656E74692E2044756973206C6967756C612066656C69732C2065666669;
        inPKT[586]      = 272'hC74A63697475722065742076656C69742061742C20666163696C6973697320636F6E;
        inPKT[587]      = 272'hC74B76616C6C6973206A7573746F2E204E756C6C616D206C6F626F72746973207065;
        inPKT[588]      = 272'hC74C6C6C656E74657371756520736F6C6C696369747564696E2E204E616D20736974;
        inPKT[589]      = 272'hC74D20616D657420646F6C6F722073697420616D6574206C656374757320696D7065;
        inPKT[590]      = 272'hC74E726469657420636F6E7365717561742E20416C697175616D206C756374757320;
        inPKT[591]      = 272'hC74F7363656C657269737175652070757275732C206964206672696E67696C6C6120;
        inPKT[592]      = 272'hC75073656D20766F6C75747061742061632E205365642074656D706F722C20656E69;
        inPKT[593]      = 272'hC7516D206567657420657569736D6F6420666163696C697369732C206E6973692065;
        inPKT[594]      = 272'hC752782073656D70657220697073756D2C20696E207361676974746973206F726369;
        inPKT[595]      = 272'hC753207175616D20696E206C65637475732E20557420766974616520656C6974206C;
        inPKT[596]      = 272'hC7546967756C612E204E756E6320656765737461732C206D69207669746165206961;
        inPKT[597]      = 272'hC75563756C6973206D61747469732C20647569206E69626820656C656966656E6420;
        inPKT[598]      = 272'hC7566E69736C2C206567657420706F727461206C696265726F206175677565207175;
        inPKT[599]      = 272'hC757697320656E696D2E205365642073697420616D65742070756C76696E61722065;
        inPKT[600]      = 272'hC758782C2076656C2070656C6C656E746573717565206C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
