`include "SIMON_defintions.svh"

module test_SIMON_4896_THROUGHPUT;

//	INPUTS
logic				clk, nR;
logic				in_newPKT;
logic				out_readPKT;
logic [(1+(`N/2)):0][7:0]	in;

//	OUTPUTS
logic 				in_loadPKT, in_donePKT;
logic				out_donePKT;
logic [(1+(`N/2)):0][7:0]	out;

SIMON_topPKT			topPKT(.*);

logic				encrypt, doneSIM;
int				countIN, countOUT, countCYCLE;

initial
begin
	#50ns		clk = 1'b0;
	forever #50ns	clk = ~clk;
end

`define				PKT_MAX 1600
logic [`PKT_MAX:0][(1+(`N/2)):0][7:0]inPKT;

initial
begin
	nR = 1'b0;	
	@(posedge clk);
	#10ns
	
	in_newPKT = 1'b0;
	out_readPKT = 1'b0;
	encrypt = 1'b1;
	doneSIM = 1'b0;
	countIN = 0;
	countOUT = 0;
	countCYCLE = 0;

        inPKT[0]        = 112'hE2001A19181211100A0908020100;
        inPKT[1]        = 112'hC2014C6F72656D20697073756D20;
        inPKT[2]        = 112'hC202646F6C6F722073697420616D;
        inPKT[3]        = 112'hC20365742C20636F6E7365637465;
        inPKT[4]        = 112'hC204747572206164697069736369;
        inPKT[5]        = 112'hC2056E6720656C69742E20437572;
        inPKT[6]        = 112'hC20661626974757220756C6C616D;
        inPKT[7]        = 112'hC207636F727065722074656D7075;
        inPKT[8]        = 112'hC20873206E6973692C2065742070;
        inPKT[9]        = 112'hC2096F73756572652075726E612E;
        inPKT[10]       = 112'hC20A2041656E65616E2073656420;
        inPKT[11]       = 112'hC20B67726176696461206C616375;
        inPKT[12]       = 112'hC20C732E204E756C6C6120666163;
        inPKT[13]       = 112'hC20D696C6973692E204E756C6C61;
        inPKT[14]       = 112'hC20E2074656D707573206F726369;
        inPKT[15]       = 112'hC20F207175697320656C69742066;
        inPKT[16]       = 112'hC2106575676961742C2076656C20;
        inPKT[17]       = 112'hC21173656D706572206C656F2069;
        inPKT[18]       = 112'hC2126D706572646965742E204D61;
        inPKT[19]       = 112'hC2136563656E6173206574206E75;
        inPKT[20]       = 112'hC2146E6320696E206E6962682066;
        inPKT[21]       = 112'hC2156163696C6973697320636F6E;
        inPKT[22]       = 112'hC21676616C6C69732E2053656420;
        inPKT[23]       = 112'hC217636F6E6775652068656E6472;
        inPKT[24]       = 112'hC2186572697420696163756C6973;
        inPKT[25]       = 112'hC2192E20566976616D7573207665;
        inPKT[26]       = 112'hC21A686963756C61206C75637475;
        inPKT[27]       = 112'hC21B73206573742C207669746165;
        inPKT[28]       = 112'hC21C207375736369706974206E69;
        inPKT[29]       = 112'hC21D736C20706F72747469746F72;
        inPKT[30]       = 112'hC21E2061632E0D0A0D0A446F6E65;
        inPKT[31]       = 112'hC21F63206D6F6C65737469652073;
        inPKT[32]       = 112'hC220617069656E2069642076756C;
        inPKT[33]       = 112'hC221707574617465207665737469;
        inPKT[34]       = 112'hC22262756C756D2E204E756C6C61;
        inPKT[35]       = 112'hC22320696E206C6967756C612066;
        inPKT[36]       = 112'hC22472696E67696C6C612C20756C;
        inPKT[37]       = 112'hC2256C616D636F72706572207572;
        inPKT[38]       = 112'hC2266E612065742C20706F727474;
        inPKT[39]       = 112'hC22769746F72206C65637475732E;
        inPKT[40]       = 112'hC228205175697371756520626C61;
        inPKT[41]       = 112'hC2296E646974206575206D617572;
        inPKT[42]       = 112'hC22A69732061632068656E647265;
        inPKT[43]       = 112'hC22B7269742E204E756C6C612076;
        inPKT[44]       = 112'hC22C656E656E617469732C206D65;
        inPKT[45]       = 112'hC22D747573206574206C75637475;
        inPKT[46]       = 112'hC22E73206672696E67696C6C612C;
        inPKT[47]       = 112'hC22F206E6962682076656C697420;
        inPKT[48]       = 112'hC230756C6C616D636F7270657220;
        inPKT[49]       = 112'hC2316469616D2C20656765742065;
        inPKT[50]       = 112'hC232666669636974757220697073;
        inPKT[51]       = 112'hC233756D20747572706973206174;
        inPKT[52]       = 112'hC234206E6962682E205574206567;
        inPKT[53]       = 112'hC2356574207072657469756D2065;
        inPKT[54]       = 112'hC236726F732C2065676574206469;
        inPKT[55]       = 112'hC2376374756D206C616375732E20;
        inPKT[56]       = 112'hC2384D616563656E617320757420;
        inPKT[57]       = 112'hC239656E696D2065782E2041656E;
        inPKT[58]       = 112'hC23A65616E207669746165207365;
        inPKT[59]       = 112'hC23B6D7065722066656C69732C20;
        inPKT[60]       = 112'hC23C73656420756C747269636965;
        inPKT[61]       = 112'hC23D732072697375732E20446F6E;
        inPKT[62]       = 112'hC23E656320636F6E736563746574;
        inPKT[63]       = 112'hC23F7572206D69206E69736C2C20;
        inPKT[64]       = 112'hC240617420637572737573206970;
        inPKT[65]       = 112'hC24173756D206772617669646120;
        inPKT[66]       = 112'hC242612E2050686173656C6C7573;
        inPKT[67]       = 112'hC2432073697420616D6574206D61;
        inPKT[68]       = 112'hC244676E612076656C2069707375;
        inPKT[69]       = 112'hC2456D206567657374617320706F;
        inPKT[70]       = 112'hC2467274612E20566976616D7573;
        inPKT[71]       = 112'hC247206C756374757320656E696D;
        inPKT[72]       = 112'hC24820656765742074656D706F72;
        inPKT[73]       = 112'hC2492073616769747469732E2041;
        inPKT[74]       = 112'hC24A6C697175616D20626962656E;
        inPKT[75]       = 112'hC24B64756D2073656D206120636F;
        inPKT[76]       = 112'hC24C6E7365637465747572206566;
        inPKT[77]       = 112'hC24D666963697475722E20446F6E;
        inPKT[78]       = 112'hC24E6563207363656C6572697371;
        inPKT[79]       = 112'hC24F756520616C697175616D2063;
        inPKT[80]       = 112'hC25075727375732E204375726162;
        inPKT[81]       = 112'hC251697475722073697420616D65;
        inPKT[82]       = 112'hC2527420626962656E64756D2065;
        inPKT[83]       = 112'hC2536C69742E2053656420646961;
        inPKT[84]       = 112'hC2546D206A7573746F2C20696163;
        inPKT[85]       = 112'hC255756C69732071756973206E75;
        inPKT[86]       = 112'hC2566C6C612076697461652C2061;
        inPKT[87]       = 112'hC2576C697175616D20657569736D;
        inPKT[88]       = 112'hC2586F642066656C69732E0D0A0D;
        inPKT[89]       = 112'hC2590A50726F696E206461706962;
        inPKT[90]       = 112'hC25A75732C206469616D2076756C;
        inPKT[91]       = 112'hC25B707574617465206672696E67;
        inPKT[92]       = 112'hC25C696C6C61206D616C65737561;
        inPKT[93]       = 112'hC25D64612C206A7573746F207075;
        inPKT[94]       = 112'hC25E72757320636F6D6D6F646F20;
        inPKT[95]       = 112'hC25F646F6C6F722C207574206469;
        inPKT[96]       = 112'hC2606374756D2065726174206E75;
        inPKT[97]       = 112'hC2616E632072757472756D207572;
        inPKT[98]       = 112'hC2626E612E204E756C6C61206772;
        inPKT[99]       = 112'hC26361766964612075726E612076;
        inPKT[100]      = 112'hC2646974616520696D7065726469;
        inPKT[101]      = 112'hC2656574206C616F726565742E20;
        inPKT[102]      = 112'hC26650656C6C656E746573717565;
        inPKT[103]      = 112'hC2672072686F6E63757320626962;
        inPKT[104]      = 112'hC268656E64756D206E6962682C20;
        inPKT[105]      = 112'hC2696964206D6F6C6C6973206469;
        inPKT[106]      = 112'hC26A616D20737573636970697420;
        inPKT[107]      = 112'hC26B61632E2050656C6C656E7465;
        inPKT[108]      = 112'hC26C737175652076656C20696163;
        inPKT[109]      = 112'hC26D756C6973206475692E204D6F;
        inPKT[110]      = 112'hC26E72626920617420616C697175;
        inPKT[111]      = 112'hC26F6574206D617373612E205072;
        inPKT[112]      = 112'hC2706F696E207669746165206F72;
        inPKT[113]      = 112'hC2716E617265206F64696F2C2065;
        inPKT[114]      = 112'hC272752076756C70757461746520;
        inPKT[115]      = 112'hC273697073756D2E2050726F696E;
        inPKT[116]      = 112'hC274206C6F626F727469732C2073;
        inPKT[117]      = 112'hC275656D206E656320657569736D;
        inPKT[118]      = 112'hC2766F642074696E636964756E74;
        inPKT[119]      = 112'hC2772C206175677565206D617572;
        inPKT[120]      = 112'hC2786973207363656C6572697371;
        inPKT[121]      = 112'hC2797565206D61676E612C206574;
        inPKT[122]      = 112'hC27A20706F7375657265206D6920;
        inPKT[123]      = 112'hC27B6E69736C206E6563206E6973;
        inPKT[124]      = 112'hC27C692E20467573636520656C69;
        inPKT[125]      = 112'hC27D74206E657175652C20766172;
        inPKT[126]      = 112'hC27E697573206574206672696E67;
        inPKT[127]      = 112'hC27F696C6C612076697461652C20;
        inPKT[128]      = 112'hC2807661726975732076656C206E;
        inPKT[129]      = 112'hC281657175652E204E756C6C6120;
        inPKT[130]      = 112'hC28265742074656D707573206A75;
        inPKT[131]      = 112'hC28373746F2E204D6F7262692075;
        inPKT[132]      = 112'hC2846C6C616D636F727065722073;
        inPKT[133]      = 112'hC2857573636970697420636F6E67;
        inPKT[134]      = 112'hC28675652E2053656420656C6569;
        inPKT[135]      = 112'hC28766656E64206F64696F206163;
        inPKT[136]      = 112'hC288207375736369706974206469;
        inPKT[137]      = 112'hC289676E697373696D2E20517569;
        inPKT[138]      = 112'hC28A7371756520616E746520656E;
        inPKT[139]      = 112'hC28B696D2C20626C616E64697420;
        inPKT[140]      = 112'hC28C696E20636F6E736571756174;
        inPKT[141]      = 112'hC28D2061632C20696E7465726475;
        inPKT[142]      = 112'hC28E6D2076697461652070757275;
        inPKT[143]      = 112'hC28F732E204D6175726973206575;
        inPKT[144]      = 112'hC29069736D6F6420706F73756572;
        inPKT[145]      = 112'hC29165206C65637475732E205669;
        inPKT[146]      = 112'hC29276616D757320696E74657264;
        inPKT[147]      = 112'hC293756D207175616D2065752073;
        inPKT[148]      = 112'hC294656D70657220666175636962;
        inPKT[149]      = 112'hC29575732E0D0A0D0A496E206D6F;
        inPKT[150]      = 112'hC2966C6573746965206E756C6C61;
        inPKT[151]      = 112'hC29720616E74652C20616320696E;
        inPKT[152]      = 112'hC29874657264756D206D61676E61;
        inPKT[153]      = 112'hC29920636F6E64696D656E74756D;
        inPKT[154]      = 112'hC29A20636F6E64696D656E74756D;
        inPKT[155]      = 112'hC29B2E204475697320756C747269;
        inPKT[156]      = 112'hC29C6369657320736F64616C6573;
        inPKT[157]      = 112'hC29D206E756C6C612C2073697420;
        inPKT[158]      = 112'hC29E616D657420756C6C616D636F;
        inPKT[159]      = 112'hC29F72706572206F64696F207072;
        inPKT[160]      = 112'hC2A0657469756D206E65632E2046;
        inPKT[161]      = 112'hC2A1757363652073656420726973;
        inPKT[162]      = 112'hC2A275732070656C6C656E746573;
        inPKT[163]      = 112'hC2A37175652C20636F6E76616C6C;
        inPKT[164]      = 112'hC2A469732073656D20656765742C;
        inPKT[165]      = 112'hC2A52068656E6472657269742065;
        inPKT[166]      = 112'hC2A67261742E204D6F7262692073;
        inPKT[167]      = 112'hC2A76F64616C6573207665686963;
        inPKT[168]      = 112'hC2A8756C61206C6F626F72746973;
        inPKT[169]      = 112'hC2A92E2041656E65616E20612074;
        inPKT[170]      = 112'hC2AA6F72746F7220637572737573;
        inPKT[171]      = 112'hC2AB2C207363656C657269737175;
        inPKT[172]      = 112'hC2AC65206C6967756C6120706F72;
        inPKT[173]      = 112'hC2AD747469746F722C2065676573;
        inPKT[174]      = 112'hC2AE7461732065726F732E204475;
        inPKT[175]      = 112'hC2AF69732074696E636964756E74;
        inPKT[176]      = 112'hC2B020746F72746F722069642070;
        inPKT[177]      = 112'hC2B16F7375657265206772617669;
        inPKT[178]      = 112'hC2B264612E20496E20636F6E7661;
        inPKT[179]      = 112'hC2B36C6C6973206D692069642069;
        inPKT[180]      = 112'hC2B47073756D206D616C65737561;
        inPKT[181]      = 112'hC2B564612C207574206469637475;
        inPKT[182]      = 112'hC2B66D2065726F7320696D706572;
        inPKT[183]      = 112'hC2B7646965742E2050726F696E20;
        inPKT[184]      = 112'hC2B8756C6C616D636F727065722C;
        inPKT[185]      = 112'hC2B9206D61757269732069642076;
        inPKT[186]      = 112'hC2BA617269757320636F6E677565;
        inPKT[187]      = 112'hC2BB2C2065726F73207361706965;
        inPKT[188]      = 112'hC2BC6E2072686F6E637573206D69;
        inPKT[189]      = 112'hC2BD2C20617420617563746F7220;
        inPKT[190]      = 112'hC2BE6E657175652061726375206C;
        inPKT[191]      = 112'hC2BF616F72656574206469616D2E;
        inPKT[192]      = 112'hC2C00D0A0D0A467573636520706F;
        inPKT[193]      = 112'hC2C172747469746F72206C696265;
        inPKT[194]      = 112'hC2C2726F20617263752C206C6163;
        inPKT[195]      = 112'hC2C3696E69612068656E64726572;
        inPKT[196]      = 112'hC2C46974206469616D20636F6E76;
        inPKT[197]      = 112'hC2C5616C6C6973207365642E2050;
        inPKT[198]      = 112'hC2C6686173656C6C7573206E6F6E;
        inPKT[199]      = 112'hC2C7207475727069732070686172;
        inPKT[200]      = 112'hC2C8657472612C20756C6C616D63;
        inPKT[201]      = 112'hC2C96F72706572206E6571756520;
        inPKT[202]      = 112'hC2CA76656C2C20736F6C6C696369;
        inPKT[203]      = 112'hC2CB747564696E2076656C69742E;
        inPKT[204]      = 112'hC2CC2050656C6C656E7465737175;
        inPKT[205]      = 112'hC2CD65206861626974616E74206D;
        inPKT[206]      = 112'hC2CE6F7262692074726973746971;
        inPKT[207]      = 112'hC2CF75652073656E656374757320;
        inPKT[208]      = 112'hC2D06574206E6574757320657420;
        inPKT[209]      = 112'hC2D16D616C657375616461206661;
        inPKT[210]      = 112'hC2D26D6573206163207475727069;
        inPKT[211]      = 112'hC2D37320656765737461732E204E;
        inPKT[212]      = 112'hC2D4616D206E6563207361706965;
        inPKT[213]      = 112'hC2D56E206D6F6C65737469652C20;
        inPKT[214]      = 112'hC2D664696374756D206D61737361;
        inPKT[215]      = 112'hC2D720656765742C206567657374;
        inPKT[216]      = 112'hC2D86173206F64696F2E20457469;
        inPKT[217]      = 112'hC2D9616D20617263752073617069;
        inPKT[218]      = 112'hC2DA656E2C207072657469756D20;
        inPKT[219]      = 112'hC2DB61206D6F6C6C697320612C20;
        inPKT[220]      = 112'hC2DC76756C707574617465206E6F;
        inPKT[221]      = 112'hC2DD6E20657261742E2055742076;
        inPKT[222]      = 112'hC2DE69746165206E696268206C6F;
        inPKT[223]      = 112'hC2DF626F72746973206C65637475;
        inPKT[224]      = 112'hC2E0732066617563696275732070;
        inPKT[225]      = 112'hC2E16F7274612065752073697420;
        inPKT[226]      = 112'hC2E2616D6574206E69736C2E204D;
        inPKT[227]      = 112'hC2E36F72626920706F7274746974;
        inPKT[228]      = 112'hC2E46F722076656C697420657520;
        inPKT[229]      = 112'hC2E5646F6C6F72206C616F726565;
        inPKT[230]      = 112'hC2E6742C2073697420616D657420;
        inPKT[231]      = 112'hC2E7696D7065726469657420656E;
        inPKT[232]      = 112'hC2E8696D20736F64616C65732E20;
        inPKT[233]      = 112'hC2E94E756C6C616D20756C6C616D;
        inPKT[234]      = 112'hC2EA636F72706572207475727069;
        inPKT[235]      = 112'hC2EB732061742070656C6C656E74;
        inPKT[236]      = 112'hC2EC657371756520766172697573;
        inPKT[237]      = 112'hC2ED2E20566976616D7573206575;
        inPKT[238]      = 112'hC2EE20696D70657264696574206E;
        inPKT[239]      = 112'hC2EF657175652E20536564207175;
        inPKT[240]      = 112'hC2F0697320617563746F7220616E;
        inPKT[241]      = 112'hC2F174652E204D61757269732073;
        inPKT[242]      = 112'hC2F2656D70657220697073756D20;
        inPKT[243]      = 112'hC2F37365642064756920706F7375;
        inPKT[244]      = 112'hC2F46572652C20617420616C6971;
        inPKT[245]      = 112'hC2F575616D206D6574757320656C;
        inPKT[246]      = 112'hC2F6656966656E642E204E756C6C;
        inPKT[247]      = 112'hC2F7616D20747269737469717565;
        inPKT[248]      = 112'hC2F820656C656966656E64206572;
        inPKT[249]      = 112'hC2F96F732C206567657420666572;
        inPKT[250]      = 112'hC2FA6D656E74756D20697073756D;
        inPKT[251]      = 112'hC2FB20656C656D656E74756D206E;
        inPKT[252]      = 112'hC2FC65632E0D0A0D0A50656C6C65;
        inPKT[253]      = 112'hC2FD6E7465737175652068656E64;
        inPKT[254]      = 112'hC2FE726572697420626962656E64;
        inPKT[255]      = 112'hC2FF756D206C6967756C612C2065;
        inPKT[256]      = 112'hC2007420736F64616C6573206D61;
        inPKT[257]      = 112'hC201676E61206461706962757320;
        inPKT[258]      = 112'hC202696E2E20496E20616C697175;
        inPKT[259]      = 112'hC203657420746F72746F72206567;
        inPKT[260]      = 112'hC204657420636F6E736563746574;
        inPKT[261]      = 112'hC205757220636F6E736563746574;
        inPKT[262]      = 112'hC20675722E205175697371756520;
        inPKT[263]      = 112'hC207747269737469717565207269;
        inPKT[264]      = 112'hC20873757320657261742C206574;
        inPKT[265]      = 112'hC20920616C697175657420656C69;
        inPKT[266]      = 112'hC20A7420616C6971756574206575;
        inPKT[267]      = 112'hC20B2E20496E7465676572206E6F;
        inPKT[268]      = 112'hC20C6E206D61676E6120696E2066;
        inPKT[269]      = 112'hC20D656C697320706F7274746974;
        inPKT[270]      = 112'hC20E6F722073616769747469732E;
        inPKT[271]      = 112'hC20F205175697371756520766976;
        inPKT[272]      = 112'hC21065727261206F726369206163;
        inPKT[273]      = 112'hC2112072757472756D206C616F72;
        inPKT[274]      = 112'hC2126565742E2041656E65616E20;
        inPKT[275]      = 112'hC213636F6E76616C6C6973206469;
        inPKT[276]      = 112'hC2146374756D207475727069732C;
        inPKT[277]      = 112'hC2152065742066696E6962757320;
        inPKT[278]      = 112'hC21673617069656E20636F6E6775;
        inPKT[279]      = 112'hC2176520696E2E20536564206120;
        inPKT[280]      = 112'hC21865726174206F726E6172652C;
        inPKT[281]      = 112'hC219206D6F6C6C6973206E69736C;
        inPKT[282]      = 112'hC21A2061632C206469676E697373;
        inPKT[283]      = 112'hC21B696D206E657175652E205175;
        inPKT[284]      = 112'hC21C6973717565206D616C657375;
        inPKT[285]      = 112'hC21D61646120706F737565726520;
        inPKT[286]      = 112'hC21E74757270697320657520756C;
        inPKT[287]      = 112'hC21F6C616D636F727065722E2044;
        inPKT[288]      = 112'hC2206F6E65632076697665727261;
        inPKT[289]      = 112'hC22120626962656E64756D206E75;
        inPKT[290]      = 112'hC2226E632C2064696374756D2069;
        inPKT[291]      = 112'hC2236D70657264696574206E6571;
        inPKT[292]      = 112'hC2247565206D6178696D75732069;
        inPKT[293]      = 112'hC2256E2E20446F6E656320757420;
        inPKT[294]      = 112'hC226756C74726963657320646F6C;
        inPKT[295]      = 112'hC2276F722E20566976616D757320;
        inPKT[296]      = 112'hC228736564206175677565207072;
        inPKT[297]      = 112'hC229657469756D2C20766F6C7574;
        inPKT[298]      = 112'hC22A70617420657261742061632C;
        inPKT[299]      = 112'hC22B20706F727461206469616D2E;
        inPKT[300]      = 112'hC22C204D617572697320696E2070;
        inPKT[301]      = 112'hC22D7572757320756C7472696369;
        inPKT[302]      = 112'hC22E65732C207375736369706974;
        inPKT[303]      = 112'hC22F206469616D207365642C2074;
        inPKT[304]      = 112'hC230696E636964756E7420656E69;
        inPKT[305]      = 112'hC2316D2E20446F6E656320717569;
        inPKT[306]      = 112'hC2327320706F7375657265206E69;
        inPKT[307]      = 112'hC23362682E20496E206861632068;
        inPKT[308]      = 112'hC234616269746173736520706C61;
        inPKT[309]      = 112'hC2357465612064696374756D7374;
        inPKT[310]      = 112'hC2362E0D0A0D0A4D6F726269206F;
        inPKT[311]      = 112'hC237726E617265206A7573746F20;
        inPKT[312]      = 112'hC2386174207175616D2066617563;
        inPKT[313]      = 112'hC239696275732C2073697420616D;
        inPKT[314]      = 112'hC23A6574206D6F6C657374696520;
        inPKT[315]      = 112'hC23B6C656F206375727375732E20;
        inPKT[316]      = 112'hC23C4D6175726973206C616F7265;
        inPKT[317]      = 112'hC23D657420616E74652061206D65;
        inPKT[318]      = 112'hC23E747573206566666963697475;
        inPKT[319]      = 112'hC23F72207661726975732E205365;
        inPKT[320]      = 112'hC240642076656C206F7263692073;
        inPKT[321]      = 112'hC24161676974746973206E756E63;
        inPKT[322]      = 112'hC24220626C616E64697420636F6E;
        inPKT[323]      = 112'hC2437365717561742E2050726165;
        inPKT[324]      = 112'hC24473656E74206D616C65737561;
        inPKT[325]      = 112'hC2456461206E6571756520717569;
        inPKT[326]      = 112'hC246732064696374756D20646967;
        inPKT[327]      = 112'hC2476E697373696D2E20446F6E65;
        inPKT[328]      = 112'hC2486320666163696C6973697320;
        inPKT[329]      = 112'hC24973697420616D65742076656C;
        inPKT[330]      = 112'hC24A6974206575206C6F626F7274;
        inPKT[331]      = 112'hC24B69732E204E756C6C616D2062;
        inPKT[332]      = 112'hC24C6C616E64697420656C656D65;
        inPKT[333]      = 112'hC24D6E74756D206D61757269732C;
        inPKT[334]      = 112'hC24E20766974616520656C656D65;
        inPKT[335]      = 112'hC24F6E74756D20646F6C6F722068;
        inPKT[336]      = 112'hC250656E64726572697420766974;
        inPKT[337]      = 112'hC25161652E204675736365206D6F;
        inPKT[338]      = 112'hC2526C65737469652C20656C6974;
        inPKT[339]      = 112'hC25320757420616C697175657420;
        inPKT[340]      = 112'hC254766F6C75747061742C206E65;
        inPKT[341]      = 112'hC2557175652076656C6974207072;
        inPKT[342]      = 112'hC256657469756D2061756775652C;
        inPKT[343]      = 112'hC257206672696E67696C6C612063;
        inPKT[344]      = 112'hC2586F6E64696D656E74756D206A;
        inPKT[345]      = 112'hC2597573746F2073617069656E20;
        inPKT[346]      = 112'hC25A61206A7573746F2E20506861;
        inPKT[347]      = 112'hC25B73656C6C7573207175697320;
        inPKT[348]      = 112'hC25C617563746F72206C6F72656D;
        inPKT[349]      = 112'hC25D2C20696E20616C697175616D;
        inPKT[350]      = 112'hC25E206E756E632E20557420656C;
        inPKT[351]      = 112'hC25F656966656E6420616E746520;
        inPKT[352]      = 112'hC2606574206E697369206D6F6C65;
        inPKT[353]      = 112'hC2617374696520636F6E76616C6C;
        inPKT[354]      = 112'hC26269732069642065742073656D;
        inPKT[355]      = 112'hC2632E2053656420616320626962;
        inPKT[356]      = 112'hC264656E64756D20617263752E20;
        inPKT[357]      = 112'hC265467573636520766573746962;
        inPKT[358]      = 112'hC266756C756D206E756E63206567;
        inPKT[359]      = 112'hC26765742074656C6C7573206665;
        inPKT[360]      = 112'hC268726D656E74756D2C206E6563;
        inPKT[361]      = 112'hC2692072686F6E637573206D6173;
        inPKT[362]      = 112'hC26A736120636F6D6D6F646F2E20;
        inPKT[363]      = 112'hC26B4D616563656E617320696420;
        inPKT[364]      = 112'hC26C6E756E63206E6F6E20657820;
        inPKT[365]      = 112'hC26D766573746962756C756D206F;
        inPKT[366]      = 112'hC26E726E617265207574206E6563;
        inPKT[367]      = 112'hC26F2065726F732E20416C697175;
        inPKT[368]      = 112'hC270616D20656666696369747572;
        inPKT[369]      = 112'hC27120636F6D6D6F646F20646961;
        inPKT[370]      = 112'hC2726D206964206C6F626F727469;
        inPKT[371]      = 112'hC273732E20536564206163207465;
        inPKT[372]      = 112'hC2746D706F72206C65637475732E;
        inPKT[373]      = 112'hC275204E756E6320656C656D656E;
        inPKT[374]      = 112'hC27674756D207574206C65637475;
        inPKT[375]      = 112'hC277732061632074696E63696475;
        inPKT[376]      = 112'hC2786E742E20557420696163756C;
        inPKT[377]      = 112'hC2796973206E756C6C6120717569;
        inPKT[378]      = 112'hC27A7320657820656C656D656E74;
        inPKT[379]      = 112'hC27B756D2C20616C697175657420;
        inPKT[380]      = 112'hC27C73656D706572206D61676E61;
        inPKT[381]      = 112'hC27D20656C656966656E642E0D0A;
        inPKT[382]      = 112'hC27E0D0A43757261626974757220;
        inPKT[383]      = 112'hC27F746F72746F72206E69736C2C;
        inPKT[384]      = 112'hC28020756C747269636965732069;
        inPKT[385]      = 112'hC2816E206E657175652061632C20;
        inPKT[386]      = 112'hC282616363756D73616E20636F6E;
        inPKT[387]      = 112'hC283736571756174206D65747573;
        inPKT[388]      = 112'hC2842E204D616563656E6173206D;
        inPKT[389]      = 112'hC285617373612073617069656E2C;
        inPKT[390]      = 112'hC286206D617474697320696E2076;
        inPKT[391]      = 112'hC287656E656E6174697320736974;
        inPKT[392]      = 112'hC28820616D65742C20617563746F;
        inPKT[393]      = 112'hC289722073697420616D65742065;
        inPKT[394]      = 112'hC28A6E696D2E204E756E63207669;
        inPKT[395]      = 112'hC28B746165206D6574757320636F;
        inPKT[396]      = 112'hC28C6D6D6F646F2C206D61747469;
        inPKT[397]      = 112'hC28D73206D617373612073697420;
        inPKT[398]      = 112'hC28E616D65742C20766172697573;
        inPKT[399]      = 112'hC28F206C6F72656D2E204E756E63;
        inPKT[400]      = 112'hC29020696E20656C697420656C69;
        inPKT[401]      = 112'hC291742E204E756E63206F726E61;
        inPKT[402]      = 112'hC292726520636F6E736563746574;
        inPKT[403]      = 112'hC2937572206D61676E612C207369;
        inPKT[404]      = 112'hC2947420616D657420706F727474;
        inPKT[405]      = 112'hC29569746F722061726375207268;
        inPKT[406]      = 112'hC2966F6E6375732065752E205375;
        inPKT[407]      = 112'hC2977370656E6469737365207363;
        inPKT[408]      = 112'hC298656C6572697371756520756C;
        inPKT[409]      = 112'hC299747269636965732065782061;
        inPKT[410]      = 112'hC29A20616C697175616D2E205375;
        inPKT[411]      = 112'hC29B7370656E6469737365207275;
        inPKT[412]      = 112'hC29C7472756D20736F6C6C696369;
        inPKT[413]      = 112'hC29D747564696E206E756E632C20;
        inPKT[414]      = 112'hC29E6E6F6E20636F6E76616C6C69;
        inPKT[415]      = 112'hC29F7320747572706973206C616F;
        inPKT[416]      = 112'hC2A0726565742073697420616D65;
        inPKT[417]      = 112'hC2A1742E2041656E65616E206120;
        inPKT[418]      = 112'hC2A266696E69627573206D617572;
        inPKT[419]      = 112'hC2A369732C207175697320637572;
        inPKT[420]      = 112'hC2A4737573206E756E632E20496E;
        inPKT[421]      = 112'hC2A5206665756769617420647569;
        inPKT[422]      = 112'hC2A62076656C2075726E61207365;
        inPKT[423]      = 112'hC2A76D7065722066617563696275;
        inPKT[424]      = 112'hC2A8732E204D617572697320756C;
        inPKT[425]      = 112'hC2A9747269636965732061742074;
        inPKT[426]      = 112'hC2AA757270697320656765742070;
        inPKT[427]      = 112'hC2AB656C6C656E7465737175652E;
        inPKT[428]      = 112'hC2AC205072616573656E74207369;
        inPKT[429]      = 112'hC2AD7420616D6574206C6967756C;
        inPKT[430]      = 112'hC2AE6120636F6E76616C6C69732C;
        inPKT[431]      = 112'hC2AF20656C656D656E74756D206E;
        inPKT[432]      = 112'hC2B0756C6C6120756C6C616D636F;
        inPKT[433]      = 112'hC2B1727065722C20616C69717561;
        inPKT[434]      = 112'hC2B26D2075726E612E2045746961;
        inPKT[435]      = 112'hC2B36D207175616D20656C69742C;
        inPKT[436]      = 112'hC2B420706F737565726520757420;
        inPKT[437]      = 112'hC2B57175616D20656765742C2066;
        inPKT[438]      = 112'hC2B6696E6962757320736F6C6C69;
        inPKT[439]      = 112'hC2B76369747564696E206E756C6C;
        inPKT[440]      = 112'hC2B8612E20496E20737573636970;
        inPKT[441]      = 112'hC2B9697420656E696D2065742065;
        inPKT[442]      = 112'hC2BA726F732066696E696275732C;
        inPKT[443]      = 112'hC2BB207574207363656C65726973;
        inPKT[444]      = 112'hC2BC7175652074656C6C75732066;
        inPKT[445]      = 112'hC2BD6575676961742E2043757261;
        inPKT[446]      = 112'hC2BE6269747572206E6F6E206D61;
        inPKT[447]      = 112'hC2BF737361207661726975732064;
        inPKT[448]      = 112'hC2C06F6C6F722067726176696461;
        inPKT[449]      = 112'hC2C120656C656D656E74756D2071;
        inPKT[450]      = 112'hC2C27569732075742066656C6973;
        inPKT[451]      = 112'hC2C32E2050686173656C6C757320;
        inPKT[452]      = 112'hC2C4657569736D6F642069707375;
        inPKT[453]      = 112'hC2C56D20656765742076656C6974;
        inPKT[454]      = 112'hC2C6206C6F626F727469732C2065;
        inPKT[455]      = 112'hC2C767657420706F727461206D61;
        inPKT[456]      = 112'hC2C8757269732074656D7075732E;
        inPKT[457]      = 112'hC2C92053656420696D7065726469;
        inPKT[458]      = 112'hC2CA657420766F6C757470617420;
        inPKT[459]      = 112'hC2CB74656C6C7573206575207469;
        inPKT[460]      = 112'hC2CC6E636964756E742E0D0A0D0A;
        inPKT[461]      = 112'hC2CD55742076656C206D69206174;
        inPKT[462]      = 112'hC2CE206D65747573206672696E67;
        inPKT[463]      = 112'hC2CF696C6C612067726176696461;
        inPKT[464]      = 112'hC2D02E205072616573656E742065;
        inPKT[465]      = 112'hC2D1726F73206E6962682C206375;
        inPKT[466]      = 112'hC2D2727375732065676573746173;
        inPKT[467]      = 112'hC2D32074696E636964756E742073;
        inPKT[468]      = 112'hC2D46F64616C65732C207363656C;
        inPKT[469]      = 112'hC2D565726973717565206E656320;
        inPKT[470]      = 112'hC2D666656C69732E20496E746567;
        inPKT[471]      = 112'hC2D7657220696D70657264696574;
        inPKT[472]      = 112'hC2D8206D616C657375616461206E;
        inPKT[473]      = 112'hC2D969736C20616C697175657420;
        inPKT[474]      = 112'hC2DA76656E656E617469732E2049;
        inPKT[475]      = 112'hC2DB6E7465676572207365642070;
        inPKT[476]      = 112'hC2DC6F72747469746F7220697073;
        inPKT[477]      = 112'hC2DD756D2E20496E746567657220;
        inPKT[478]      = 112'hC2DE636F6D6D6F646F2066657567;
        inPKT[479]      = 112'hC2DF69617420746F72746F722C20;
        inPKT[480]      = 112'hC2E06575206C6F626F7274697320;
        inPKT[481]      = 112'hC2E1617567756520656C656D656E;
        inPKT[482]      = 112'hC2E274756D2073697420616D6574;
        inPKT[483]      = 112'hC2E32E20446F6E65632076657374;
        inPKT[484]      = 112'hC2E46962756C756D206C6967756C;
        inPKT[485]      = 112'hC2E5612061756775652C20657420;
        inPKT[486]      = 112'hC2E666696E696275732061726375;
        inPKT[487]      = 112'hC2E720706F72746120696E2E204E;
        inPKT[488]      = 112'hC2E8756C6C612073656D2074656C;
        inPKT[489]      = 112'hC2E96C75732C20756C6C616D636F;
        inPKT[490]      = 112'hC2EA727065722061742063757273;
        inPKT[491]      = 112'hC2EB757320612C20706F72746120;
        inPKT[492]      = 112'hC2EC73697420616D6574206D6167;
        inPKT[493]      = 112'hC2ED6E612E204E756E6320766974;
        inPKT[494]      = 112'hC2EE616520696D70657264696574;
        inPKT[495]      = 112'hC2EF2070757275732C206E656320;
        inPKT[496]      = 112'hC2F0736F6C6C696369747564696E;
        inPKT[497]      = 112'hC2F12074656C6C75732E20416C69;
        inPKT[498]      = 112'hC2F27175616D206572617420766F;
        inPKT[499]      = 112'hC2F36C75747061742E2053656420;
        inPKT[500]      = 112'hC2F46964206D61676E6120636F6D;
        inPKT[501]      = 112'hC2F56D6F646F2C206C7563747573;
        inPKT[502]      = 112'hC2F62076656C697420717569732C;
        inPKT[503]      = 112'hC2F720657569736D6F6420656E69;
        inPKT[504]      = 112'hC2F86D2E20496E7465676572206D;
        inPKT[505]      = 112'hC2F9617474697320736F64616C65;
        inPKT[506]      = 112'hC2FA73206665726D656E74756D2E;
        inPKT[507]      = 112'hC2FB205175697371756520736564;
        inPKT[508]      = 112'hC2FC206672696E67696C6C61206C;
        inPKT[509]      = 112'hC2FD6F72656D2E20437261732076;
        inPKT[510]      = 112'hC2FE65686963756C612074656D70;
        inPKT[511]      = 112'hC2FF75732073617069656E207574;
        inPKT[512]      = 112'hC20020636F6E6775652E20447569;
        inPKT[513]      = 112'hC201732073617069656E20656E69;
        inPKT[514]      = 112'hC2026D2C20706F727461206E6563;
        inPKT[515]      = 112'hC203206C656F2069642C20656666;
        inPKT[516]      = 112'hC20469636974757220706F737565;
        inPKT[517]      = 112'hC2057265206C696265726F2E204E;
        inPKT[518]      = 112'hC206756C6C616D2061632074656D;
        inPKT[519]      = 112'hC207706F72206D657475732E2053;
        inPKT[520]      = 112'hC20865642076656C207475727069;
        inPKT[521]      = 112'hC2097320666575676961742C2069;
        inPKT[522]      = 112'hC20A6163756C6973206175677565;
        inPKT[523]      = 112'hC20B20717569732C2074696E6369;
        inPKT[524]      = 112'hC20C64756E74207475727069732E;
        inPKT[525]      = 112'hC20D0D0A0D0A566976616D757320;
        inPKT[526]      = 112'hC20E706F737565726520706F7274;
        inPKT[527]      = 112'hC20F7469746F722061756775652C;
        inPKT[528]      = 112'hC210207661726975732061636375;
        inPKT[529]      = 112'hC2116D73616E20656C6974207675;
        inPKT[530]      = 112'hC2126C7075746174652065676574;
        inPKT[531]      = 112'hC2132E2051756973717565207365;
        inPKT[532]      = 112'hC21464206D616C65737561646120;
        inPKT[533]      = 112'hC2156E69736C2E20496E74657264;
        inPKT[534]      = 112'hC216756D206574206D616C657375;
        inPKT[535]      = 112'hC2176164612066616D6573206163;
        inPKT[536]      = 112'hC21820616E746520697073756D20;
        inPKT[537]      = 112'hC2197072696D697320696E206661;
        inPKT[538]      = 112'hC21A7563696275732E204E756E63;
        inPKT[539]      = 112'hC21B20747572706973206469616D;
        inPKT[540]      = 112'hC21C2C2073757363697069742061;
        inPKT[541]      = 112'hC21D632065726F732076656C2C20;
        inPKT[542]      = 112'hC21E74656D7075732076656E656E;
        inPKT[543]      = 112'hC21F6174697320697073756D2E20;
        inPKT[544]      = 112'hC22044756973206C756374757320;
        inPKT[545]      = 112'hC22172686F6E637573206D617373;
        inPKT[546]      = 112'hC222612E20467573636520757420;
        inPKT[547]      = 112'hC2236C6163696E69612074757270;
        inPKT[548]      = 112'hC22469732E20566976616D757320;
        inPKT[549]      = 112'hC22572757472756D2074656C6C75;
        inPKT[550]      = 112'hC226732061756775652C20617420;
        inPKT[551]      = 112'hC2276F726E617265206E69736C20;
        inPKT[552]      = 112'hC228666163696C69736973206574;
        inPKT[553]      = 112'hC2292E204E756E6320736564206E;
        inPKT[554]      = 112'hC22A6973692072697375732E2049;
        inPKT[555]      = 112'hC22B6E746567657220656C656D65;
        inPKT[556]      = 112'hC22C6E74756D206D617572697320;
        inPKT[557]      = 112'hC22D7175616D2C20757420766568;
        inPKT[558]      = 112'hC22E6963756C61206D6175726973;
        inPKT[559]      = 112'hC22F20636F6E6775652065752E0D;
        inPKT[560]      = 112'hC2300A0D0A467573636520612074;
        inPKT[561]      = 112'hC231656C6C75732073697420616D;
        inPKT[562]      = 112'hC23265742065726174206665726D;
        inPKT[563]      = 112'hC233656E74756D207363656C6572;
        inPKT[564]      = 112'hC23469737175652E204375726162;
        inPKT[565]      = 112'hC2356974757220696E2076656C69;
        inPKT[566]      = 112'hC2367420617420656E696D206C61;
        inPKT[567]      = 112'hC23763696E696120766568696375;
        inPKT[568]      = 112'hC2386C61206163206964206A7573;
        inPKT[569]      = 112'hC239746F2E2050726F696E206E6F;
        inPKT[570]      = 112'hC23A6E20646F6C6F722065666669;
        inPKT[571]      = 112'hC23B63697475722C2074696E6369;
        inPKT[572]      = 112'hC23C64756E74206F64696F206575;
        inPKT[573]      = 112'hC23D2C2066617563696275732065;
        inPKT[574]      = 112'hC23E6E696D2E2050656C6C656E74;
        inPKT[575]      = 112'hC23F657371756520646170696275;
        inPKT[576]      = 112'hC24073206F726369206163206C6F;
        inPKT[577]      = 112'hC24172656D20696163756C69732C;
        inPKT[578]      = 112'hC2422073697420616D657420626C;
        inPKT[579]      = 112'hC243616E64697420617263752074;
        inPKT[580]      = 112'hC24472697374697175652E204165;
        inPKT[581]      = 112'hC2456E65616E2074726973746971;
        inPKT[582]      = 112'hC246756520746F72746F72206E65;
        inPKT[583]      = 112'hC24763206A7573746F20616C6971;
        inPKT[584]      = 112'hC24875616D2C20696E2070726574;
        inPKT[585]      = 112'hC24969756D2066656C6973206D6F;
        inPKT[586]      = 112'hC24A6C65737469652E2053656420;
        inPKT[587]      = 112'hC24B65742074656D707573206175;
        inPKT[588]      = 112'hC24C6775652E204E756C6C612066;
        inPKT[589]      = 112'hC24D72696E67696C6C6120656C65;
        inPKT[590]      = 112'hC24E6966656E6420697073756D20;
        inPKT[591]      = 112'hC24F766976657272612063757273;
        inPKT[592]      = 112'hC25075732E20416C697175616D20;
        inPKT[593]      = 112'hC2516D6178696D7573206665726D;
        inPKT[594]      = 112'hC252656E74756D206E6962682061;
        inPKT[595]      = 112'hC2536320616363756D73616E2E20;
        inPKT[596]      = 112'hC2544E756C6C6120666163696C69;
        inPKT[597]      = 112'hC25573692E20566573746962756C;
        inPKT[598]      = 112'hC256756D20666163696C69736973;
        inPKT[599]      = 112'hC257206C656F2065676573746173;
        inPKT[600]      = 112'hC2582073656D206D617474697320;
        inPKT[601]      = 112'hC259636F6E6775652E204D617572;
        inPKT[602]      = 112'hC25A697320766974616520657820;
        inPKT[603]      = 112'hC25B617420726973757320646170;
        inPKT[604]      = 112'hC25C6962757320656C656966656E;
        inPKT[605]      = 112'hC25D642E20496E74656765722075;
        inPKT[606]      = 112'hC25E742065726F7320636F6E6775;
        inPKT[607]      = 112'hC25F652C20706F72747469746F72;
        inPKT[608]      = 112'hC26020616E7465206E6F6E2C2069;
        inPKT[609]      = 112'hC2616E74657264756D20646F6C6F;
        inPKT[610]      = 112'hC262722E0D0A0D0A566573746962;
        inPKT[611]      = 112'hC263756C756D20656C656966656E;
        inPKT[612]      = 112'hC26464206D617572697320657520;
        inPKT[613]      = 112'hC2656E6973692064696374756D20;
        inPKT[614]      = 112'hC266677261766964612E20447569;
        inPKT[615]      = 112'hC26773206D6F6C6C697320646961;
        inPKT[616]      = 112'hC2686D2076656C20656E696D2074;
        inPKT[617]      = 112'hC269656D7075732C207669746165;
        inPKT[618]      = 112'hC26A2064617069627573206D6173;
        inPKT[619]      = 112'hC26B73612073616769747469732E;
        inPKT[620]      = 112'hC26C204E756C6C61207574206175;
        inPKT[621]      = 112'hC26D63746F7220746F72746F722E;
        inPKT[622]      = 112'hC26E204D6F72626920736564206C;
        inPKT[623]      = 112'hC26F6F72656D2075726E612E2046;
        inPKT[624]      = 112'hC27075736365206D61747469732C;
        inPKT[625]      = 112'hC271206D61676E6120616320636F;
        inPKT[626]      = 112'hC2726E64696D656E74756D206665;
        inPKT[627]      = 112'hC27375676961742C206D61737361;
        inPKT[628]      = 112'hC27420647569206D6178696D7573;
        inPKT[629]      = 112'hC275206E756C6C612C2065752061;
        inPKT[630]      = 112'hC2766C6971756574206E65717565;
        inPKT[631]      = 112'hC277206D61757269732061206572;
        inPKT[632]      = 112'hC27861742E205175697371756520;
        inPKT[633]      = 112'hC279617563746F72206573742075;
        inPKT[634]      = 112'hC27A7420696E74657264756D2063;
        inPKT[635]      = 112'hC27B6F6E73656374657475722E20;
        inPKT[636]      = 112'hC27C446F6E656320656765742064;
        inPKT[637]      = 112'hC27D69676E697373696D20746F72;
        inPKT[638]      = 112'hC27E746F722C2068656E64726572;
        inPKT[639]      = 112'hC27F6974206D6174746973206572;
        inPKT[640]      = 112'hC28061742E2050656C6C656E7465;
        inPKT[641]      = 112'hC28173717565206861626974616E;
        inPKT[642]      = 112'hC28274206D6F7262692074726973;
        inPKT[643]      = 112'hC28374697175652073656E656374;
        inPKT[644]      = 112'hC2847573206574206E6574757320;
        inPKT[645]      = 112'hC2856574206D616C657375616461;
        inPKT[646]      = 112'hC2862066616D6573206163207475;
        inPKT[647]      = 112'hC287727069732065676573746173;
        inPKT[648]      = 112'hC2882E2051756973717565206F72;
        inPKT[649]      = 112'hC2896E6172652076617269757320;
        inPKT[650]      = 112'hC28A74656D7075732E0D0A0D0A4D;
        inPKT[651]      = 112'hC28B6F7262692072757472756D20;
        inPKT[652]      = 112'hC28C616E7465206E6962682C2061;
        inPKT[653]      = 112'hC28D2076697665727261206E756C;
        inPKT[654]      = 112'hC28E6C612068656E647265726974;
        inPKT[655]      = 112'hC28F20696E2E2050726F696E2073;
        inPKT[656]      = 112'hC290757363697069742065676573;
        inPKT[657]      = 112'hC29174617320657261742C207574;
        inPKT[658]      = 112'hC29220617563746F72206F726369;
        inPKT[659]      = 112'hC293206D617474697320612E2050;
        inPKT[660]      = 112'hC294656C6C656E74657371756520;
        inPKT[661]      = 112'hC2956C7563747573206672696E67;
        inPKT[662]      = 112'hC296696C6C6120656C6974207574;
        inPKT[663]      = 112'hC297206C6163696E69612E205574;
        inPKT[664]      = 112'hC298206574206D61737361206E75;
        inPKT[665]      = 112'hC2996C6C612E2053656420617420;
        inPKT[666]      = 112'hC29A6672696E67696C6C61206C6F;
        inPKT[667]      = 112'hC29B72656D2E2050726F696E2067;
        inPKT[668]      = 112'hC29C72617669646120616363756D;
        inPKT[669]      = 112'hC29D73616E207269737573207365;
        inPKT[670]      = 112'hC29E6420626962656E64756D2E20;
        inPKT[671]      = 112'hC29F4D616563656E6173206D616C;
        inPKT[672]      = 112'hC2A0657375616461206F64696F20;
        inPKT[673]      = 112'hC2A175742076656C697420657569;
        inPKT[674]      = 112'hC2A2736D6F642064617069627573;
        inPKT[675]      = 112'hC2A32E0D0A0D0A457469616D2063;
        inPKT[676]      = 112'hC2A46F6E677565206D6174746973;
        inPKT[677]      = 112'hC2A520696163756C69732E204D61;
        inPKT[678]      = 112'hC2A6757269732076697461652065;
        inPKT[679]      = 112'hC2A766666963697475722073656D;
        inPKT[680]      = 112'hC2A82E205365642070756C76696E;
        inPKT[681]      = 112'hC2A9617220646F6C6F7220757420;
        inPKT[682]      = 112'hC2AA6D6920657569736D6F642068;
        inPKT[683]      = 112'hC2AB656E6472657269742E204E75;
        inPKT[684]      = 112'hC2AC6C6C616D2061742067726176;
        inPKT[685]      = 112'hC2AD69646120646F6C6F722E204D;
        inPKT[686]      = 112'hC2AE6F726269206C656F20747572;
        inPKT[687]      = 112'hC2AF7069732C20636F6E67756520;
        inPKT[688]      = 112'hC2B06E656320616C697175616D20;
        inPKT[689]      = 112'hC2B175742C20636F6D6D6F646F20;
        inPKT[690]      = 112'hC2B2696E206E756E632E204E756C;
        inPKT[691]      = 112'hC2B36C6120617420666175636962;
        inPKT[692]      = 112'hC2B47573206C656F2C2065752066;
        inPKT[693]      = 112'hC2B5657567696174206C61637573;
        inPKT[694]      = 112'hC2B62E204675736365206E6F6E20;
        inPKT[695]      = 112'hC2B7656765737461732074757270;
        inPKT[696]      = 112'hC2B869732E205175697371756520;
        inPKT[697]      = 112'hC2B9766974616520697073756D20;
        inPKT[698]      = 112'hC2BA6D692E204E756E63206E6F6E;
        inPKT[699]      = 112'hC2BB206F7263692073697420616D;
        inPKT[700]      = 112'hC2BC6574206E6973692076617269;
        inPKT[701]      = 112'hC2BD757320706F72747469746F72;
        inPKT[702]      = 112'hC2BE20696E2076756C7075746174;
        inPKT[703]      = 112'hC2BF6520746F72746F722E204E75;
        inPKT[704]      = 112'hC2C06E6320636F6E76616C6C6973;
        inPKT[705]      = 112'hC2C1206772617669646120646961;
        inPKT[706]      = 112'hC2C26D206120756C747269636965;
        inPKT[707]      = 112'hC2C3732E20517569737175652065;
        inPKT[708]      = 112'hC2C475206A7573746F20636F6E64;
        inPKT[709]      = 112'hC2C5696D656E74756D2C20766172;
        inPKT[710]      = 112'hC2C6697573206469616D2076656C;
        inPKT[711]      = 112'hC2C72C20766573746962756C756D;
        inPKT[712]      = 112'hC2C8206D617373612E0D0A0D0A50;
        inPKT[713]      = 112'hC2C9656C6C656E74657371756520;
        inPKT[714]      = 112'hC2CA70656C6C656E746573717565;
        inPKT[715]      = 112'hC2CB2073617069656E206E657175;
        inPKT[716]      = 112'hC2CC652C20617563746F72206D61;
        inPKT[717]      = 112'hC2CD6C6573756164612065726174;
        inPKT[718]      = 112'hC2CE2068656E647265726974206E;
        inPKT[719]      = 112'hC2CF65632E204E756C6C6120706C;
        inPKT[720]      = 112'hC2D0616365726174206469616D20;
        inPKT[721]      = 112'hC2D168656E647265726974206D61;
        inPKT[722]      = 112'hC2D273736120626962656E64756D;
        inPKT[723]      = 112'hC2D32C2061206D6F6C6573746965;
        inPKT[724]      = 112'hC2D42066656C69732068656E6472;
        inPKT[725]      = 112'hC2D5657269742E204D6175726973;
        inPKT[726]      = 112'hC2D620657569736D6F642076656E;
        inPKT[727]      = 112'hC2D7656E61746973206A7573746F;
        inPKT[728]      = 112'hC2D82C20757420617563746F7220;
        inPKT[729]      = 112'hC2D9656C697420616C6971756574;
        inPKT[730]      = 112'hC2DA2075742E2046757363652061;
        inPKT[731]      = 112'hC2DB6C69717565742C207175616D;
        inPKT[732]      = 112'hC2DC207574206469676E69737369;
        inPKT[733]      = 112'hC2DD6D2068656E6472657269742C;
        inPKT[734]      = 112'hC2DE206D61757269732074757270;
        inPKT[735]      = 112'hC2DF6973206469676E697373696D;
        inPKT[736]      = 112'hC2E020746F72746F722C20656765;
        inPKT[737]      = 112'hC2E1742070656C6C656E74657371;
        inPKT[738]      = 112'hC2E275652076656C6974206F7263;
        inPKT[739]      = 112'hC2E369206E6563207175616D2E20;
        inPKT[740]      = 112'hC2E44E756E632065676573746173;
        inPKT[741]      = 112'hC2E52070656C6C656E7465737175;
        inPKT[742]      = 112'hC2E6652072697375732E20437572;
        inPKT[743]      = 112'hC2E7616269747572207375736369;
        inPKT[744]      = 112'hC2E87069742074656D707573206C;
        inPKT[745]      = 112'hC2E9616375732C20656765742070;
        inPKT[746]      = 112'hC2EA72657469756D20656C697420;
        inPKT[747]      = 112'hC2EB74696E636964756E74206E6F;
        inPKT[748]      = 112'hC2EC6E2E20437261732075726E61;
        inPKT[749]      = 112'hC2ED206C6F72656D2C20706C6163;
        inPKT[750]      = 112'hC2EE6572617420766F6C75747061;
        inPKT[751]      = 112'hC2EF7420696D7065726469657420;
        inPKT[752]      = 112'hC2F073697420616D65742C206567;
        inPKT[753]      = 112'hC2F165737461732076656C206F72;
        inPKT[754]      = 112'hC2F263692E0D0A0D0A50656C6C65;
        inPKT[755]      = 112'hC2F36E74657371756520736F6461;
        inPKT[756]      = 112'hC2F46C6573206665726D656E7475;
        inPKT[757]      = 112'hC2F56D206E69736C2C2061742066;
        inPKT[758]      = 112'hC2F672696E67696C6C6120647569;
        inPKT[759]      = 112'hC2F72073656D706572206665726D;
        inPKT[760]      = 112'hC2F8656E74756D2E204E756C6C61;
        inPKT[761]      = 112'hC2F96D20706C6163657261742076;
        inPKT[762]      = 112'hC2FA656C206D692068656E647265;
        inPKT[763]      = 112'hC2FB72697420656C656D656E7475;
        inPKT[764]      = 112'hC2FC6D2E20457469616D206E6F6E;
        inPKT[765]      = 112'hC2FD20697073756D2065782E204E;
        inPKT[766]      = 112'hC2FE616D206163207363656C6572;
        inPKT[767]      = 112'hC2FF6973717565206E6962682C20;
        inPKT[768]      = 112'hC20076656C20666163696C697369;
        inPKT[769]      = 112'hC20173206D692E20446F6E656320;
        inPKT[770]      = 112'hC20265676573746173206C616F72;
        inPKT[771]      = 112'hC2036565742065726F732C206567;
        inPKT[772]      = 112'hC204657420766F6C757470617420;
        inPKT[773]      = 112'hC2056D657475732E205072616573;
        inPKT[774]      = 112'hC206656E7420616363756D73616E;
        inPKT[775]      = 112'hC20720626962656E64756D206E69;
        inPKT[776]      = 112'hC208736C206E65632076656E656E;
        inPKT[777]      = 112'hC209617469732E20536564207275;
        inPKT[778]      = 112'hC20A7472756D206D692061207375;
        inPKT[779]      = 112'hC20B736369706974207068617265;
        inPKT[780]      = 112'hC20C7472612E2053656420736974;
        inPKT[781]      = 112'hC20D20616D657420696E74657264;
        inPKT[782]      = 112'hC20E756D207475727069732E2041;
        inPKT[783]      = 112'hC20F6C697175616D206575206E69;
        inPKT[784]      = 112'hC210626820746F72746F722E2044;
        inPKT[785]      = 112'hC2116F6E65632066617563696275;
        inPKT[786]      = 112'hC212732064617069627573206E69;
        inPKT[787]      = 112'hC21373692C20736564206C616F72;
        inPKT[788]      = 112'hC214656574206F72636920736365;
        inPKT[789]      = 112'hC2156C6572697371756520696E2E;
        inPKT[790]      = 112'hC2160D0A0D0A4D61757269732069;
        inPKT[791]      = 112'hC2176E2066656C6973206665726D;
        inPKT[792]      = 112'hC218656E74756D2C20636F6E7661;
        inPKT[793]      = 112'hC2196C6C69732061756775652076;
        inPKT[794]      = 112'hC21A656C2C20706F737565726520;
        inPKT[795]      = 112'hC21B6D692E2050656C6C656E7465;
        inPKT[796]      = 112'hC21C73717565207363656C657269;
        inPKT[797]      = 112'hC21D737175652072686F6E637573;
        inPKT[798]      = 112'hC21E206A7573746F2C2065752070;
        inPKT[799]      = 112'hC21F756C76696E617220656E696D;
        inPKT[800]      = 112'hC2202070756C76696E6172207665;
        inPKT[801]      = 112'hC2216C2E204D616563656E617320;
        inPKT[802]      = 112'hC2227068617265747261206C6962;
        inPKT[803]      = 112'hC22365726F206D61676E612C2061;
        inPKT[804]      = 112'hC2246320736F6C6C696369747564;
        inPKT[805]      = 112'hC225696E206C656F206D6F6C6C69;
        inPKT[806]      = 112'hC22673206E6F6E2E204E756C6C61;
        inPKT[807]      = 112'hC22720656C656D656E74756D206F;
        inPKT[808]      = 112'hC228726E61726520656765737461;
        inPKT[809]      = 112'hC229732E20436C61737320617074;
        inPKT[810]      = 112'hC22A656E74207461636974692073;
        inPKT[811]      = 112'hC22B6F63696F737175206164206C;
        inPKT[812]      = 112'hC22C69746F726120746F72717565;
        inPKT[813]      = 112'hC22D6E742070657220636F6E7562;
        inPKT[814]      = 112'hC22E6961206E6F737472612C2070;
        inPKT[815]      = 112'hC22F657220696E636570746F7320;
        inPKT[816]      = 112'hC23068696D656E61656F732E2050;
        inPKT[817]      = 112'hC23172616573656E742061756775;
        inPKT[818]      = 112'hC23265206D61757269732C207268;
        inPKT[819]      = 112'hC2336F6E63757320717569732065;
        inPKT[820]      = 112'hC2347374206E6F6E2C206D6F6C6C;
        inPKT[821]      = 112'hC235697320636F6E76616C6C6973;
        inPKT[822]      = 112'hC2362066656C69732E2053757370;
        inPKT[823]      = 112'hC237656E64697373652066616369;
        inPKT[824]      = 112'hC2386C697369732C206F72636920;
        inPKT[825]      = 112'hC2397669746165206C6163696E69;
        inPKT[826]      = 112'hC23A612074656D706F722C206C65;
        inPKT[827]      = 112'hC23B637475732073617069656E20;
        inPKT[828]      = 112'hC23C6D6174746973207269737573;
        inPKT[829]      = 112'hC23D2C206E6F6E20736167697474;
        inPKT[830]      = 112'hC23E697320656C6974206E657175;
        inPKT[831]      = 112'hC23F652071756973206A7573746F;
        inPKT[832]      = 112'hC2402E20446F6E6563206D616C65;
        inPKT[833]      = 112'hC2417375616461206C6163696E69;
        inPKT[834]      = 112'hC24261206475692E205068617365;
        inPKT[835]      = 112'hC2436C6C75732068656E64726572;
        inPKT[836]      = 112'hC2446974206D6175726973206D61;
        inPKT[837]      = 112'hC245757269732C20736564206672;
        inPKT[838]      = 112'hC246696E67696C6C61206C696265;
        inPKT[839]      = 112'hC247726F206672696E67696C6C61;
        inPKT[840]      = 112'hC24820696E2E2053656420617420;
        inPKT[841]      = 112'hC2496C6967756C6120696E206A75;
        inPKT[842]      = 112'hC24A73746F2066696E6962757320;
        inPKT[843]      = 112'hC24B76756C7075746174652E204E;
        inPKT[844]      = 112'hC24C756E6320637572737573206E;
        inPKT[845]      = 112'hC24D657175652073697420616D65;
        inPKT[846]      = 112'hC24E7420617263752074696E6369;
        inPKT[847]      = 112'hC24F64756E742C20766974616520;
        inPKT[848]      = 112'hC25070686172657472612073656D;
        inPKT[849]      = 112'hC25120706F72747469746F722E20;
        inPKT[850]      = 112'hC252416C697175616D206D617474;
        inPKT[851]      = 112'hC25369732C206A7573746F206E6F;
        inPKT[852]      = 112'hC2546E20657569736D6F6420636F;
        inPKT[853]      = 112'hC2556E76616C6C69732C206E756E;
        inPKT[854]      = 112'hC25663206D6920636F6E73657175;
        inPKT[855]      = 112'hC2576174206573742C206E656320;
        inPKT[856]      = 112'hC258736F6C6C696369747564696E;
        inPKT[857]      = 112'hC259206C65637475732073617069;
        inPKT[858]      = 112'hC25A656E2076656C206F64696F2E;
        inPKT[859]      = 112'hC25B20496E2074656D706F722065;
        inPKT[860]      = 112'hC25C72617420646F6C6F722C2073;
        inPKT[861]      = 112'hC25D6564207665686963756C6120;
        inPKT[862]      = 112'hC25E75726E6120636F6E73657175;
        inPKT[863]      = 112'hC25F6174207365642E0D0A0D0A4E;
        inPKT[864]      = 112'hC260616D2072686F6E6375732069;
        inPKT[865]      = 112'hC26164206D6175726973206E6563;
        inPKT[866]      = 112'hC262206469676E697373696D2E20;
        inPKT[867]      = 112'hC263496E20696D70657264696574;
        inPKT[868]      = 112'hC26420756C747269636573206572;
        inPKT[869]      = 112'hC2656174206E656320736F6C6C69;
        inPKT[870]      = 112'hC2666369747564696E2E20496E74;
        inPKT[871]      = 112'hC267656765722073656420636F6E;
        inPKT[872]      = 112'hC26864696D656E74756D2065726F;
        inPKT[873]      = 112'hC269732E20446F6E656320656765;
        inPKT[874]      = 112'hC26A74206E756E63206964206D61;
        inPKT[875]      = 112'hC26B757269732074726973746971;
        inPKT[876]      = 112'hC26C756520706F72747469746F72;
        inPKT[877]      = 112'hC26D206C616F7265657420766974;
        inPKT[878]      = 112'hC26E6165206D657475732E204E75;
        inPKT[879]      = 112'hC26F6C6C6120666163696C697369;
        inPKT[880]      = 112'hC2702E204E756C6C616D20657520;
        inPKT[881]      = 112'hC2716C616375732061206469616D;
        inPKT[882]      = 112'hC272207472697374697175652065;
        inPKT[883]      = 112'hC273676573746173206E6F6E2069;
        inPKT[884]      = 112'hC2746163756C6973206D65747573;
        inPKT[885]      = 112'hC2752E20416C697175616D20696E;
        inPKT[886]      = 112'hC2762074656D706F722065726174;
        inPKT[887]      = 112'hC2772C20696420636F6E67756520;
        inPKT[888]      = 112'hC2786D617373612E20566976616D;
        inPKT[889]      = 112'hC27975732076656C20746F72746F;
        inPKT[890]      = 112'hC27A72207669746165206E696268;
        inPKT[891]      = 112'hC27B20636F6D6D6F646F206C6F62;
        inPKT[892]      = 112'hC27C6F7274697320717569732061;
        inPKT[893]      = 112'hC27D20697073756D2E2050726F69;
        inPKT[894]      = 112'hC27E6E20766F6C75747061742071;
        inPKT[895]      = 112'hC27F75616D206E6F6E2066656C69;
        inPKT[896]      = 112'hC280732074656D7075732C206964;
        inPKT[897]      = 112'hC28120706F737565726520646F6C;
        inPKT[898]      = 112'hC2826F722074656D706F722E2050;
        inPKT[899]      = 112'hC28372616573656E742076697461;
        inPKT[900]      = 112'hC284652074696E636964756E7420;
        inPKT[901]      = 112'hC28573617069656E2E204D616563;
        inPKT[902]      = 112'hC286656E617320666163696C6973;
        inPKT[903]      = 112'hC2876973206D617474697320616E;
        inPKT[904]      = 112'hC288746520717569732076617269;
        inPKT[905]      = 112'hC28975732E20446F6E6563207065;
        inPKT[906]      = 112'hC28A6C6C656E7465737175652065;
        inPKT[907]      = 112'hC28B726F73206665756769617420;
        inPKT[908]      = 112'hC28C74696E636964756E7420636F;
        inPKT[909]      = 112'hC28D6E64696D656E74756D2E2050;
        inPKT[910]      = 112'hC28E726F696E2066617563696275;
        inPKT[911]      = 112'hC28F7320766F6C7574706174206D;
        inPKT[912]      = 112'hC290692073656420736167697474;
        inPKT[913]      = 112'hC29169732E0D0A0D0A4475697320;
        inPKT[914]      = 112'hC2926772617669646120656C656D;
        inPKT[915]      = 112'hC293656E74756D20696E74657264;
        inPKT[916]      = 112'hC294756D2E2050726F696E207369;
        inPKT[917]      = 112'hC2957420616D6574207175616D20;
        inPKT[918]      = 112'hC2966C6967756C612E2050686173;
        inPKT[919]      = 112'hC297656C6C757320636F6D6D6F64;
        inPKT[920]      = 112'hC2986F2C2075726E6120696E2063;
        inPKT[921]      = 112'hC2996F6E67756520766F6C757470;
        inPKT[922]      = 112'hC29A61742C206C6967756C612065;
        inPKT[923]      = 112'hC29B78207068617265747261206C;
        inPKT[924]      = 112'hC29C6967756C612C20696E206469;
        inPKT[925]      = 112'hC29D6374756D206D61676E61206F;
        inPKT[926]      = 112'hC29E726369206E6563206D617572;
        inPKT[927]      = 112'hC29F69732E204E756E6320617563;
        inPKT[928]      = 112'hC2A0746F7220636F6E7365637465;
        inPKT[929]      = 112'hC2A174757220766F6C7574706174;
        inPKT[930]      = 112'hC2A22E204D6F7262692074696E63;
        inPKT[931]      = 112'hC2A36964756E74206E6962682075;
        inPKT[932]      = 112'hC2A47420656E696D206566666963;
        inPKT[933]      = 112'hC2A5697475722067726176696461;
        inPKT[934]      = 112'hC2A62E2043757261626974757220;
        inPKT[935]      = 112'hC2A77669746165207175616D2065;
        inPKT[936]      = 112'hC2A8726F732E2044756973206672;
        inPKT[937]      = 112'hC2A9696E67696C6C612061632074;
        inPKT[938]      = 112'hC2AA6F72746F7220696E2074696E;
        inPKT[939]      = 112'hC2AB636964756E742E204E756E63;
        inPKT[940]      = 112'hC2AC2076656C206D617572697320;
        inPKT[941]      = 112'hC2AD72697375732E20446F6E6563;
        inPKT[942]      = 112'hC2AE20656C656966656E64206C69;
        inPKT[943]      = 112'hC2AF67756C612073616769747469;
        inPKT[944]      = 112'hC2B073206E6973692066696E6962;
        inPKT[945]      = 112'hC2B175732C2061207363656C6572;
        inPKT[946]      = 112'hC2B26973717565206C696265726F;
        inPKT[947]      = 112'hC2B32070656C6C656E7465737175;
        inPKT[948]      = 112'hC2B4652E20566573746962756C75;
        inPKT[949]      = 112'hC2B56D2074726973746971756520;
        inPKT[950]      = 112'hC2B66D61737361206E6962682C20;
        inPKT[951]      = 112'hC2B7617420766573746962756C75;
        inPKT[952]      = 112'hC2B86D206D61676E612066696E69;
        inPKT[953]      = 112'hC2B96275732065752E0D0A0D0A43;
        inPKT[954]      = 112'hC2BA757261626974757220696D70;
        inPKT[955]      = 112'hC2BB657264696574207075727573;
        inPKT[956]      = 112'hC2BC2065676574206E756E632075;
        inPKT[957]      = 112'hC2BD6C7472696365732C20766974;
        inPKT[958]      = 112'hC2BE61652076656E656E61746973;
        inPKT[959]      = 112'hC2BF206D6173736120636F6D6D6F;
        inPKT[960]      = 112'hC2C0646F2E2050656C6C656E7465;
        inPKT[961]      = 112'hC2C173717565206861626974616E;
        inPKT[962]      = 112'hC2C274206D6F7262692074726973;
        inPKT[963]      = 112'hC2C374697175652073656E656374;
        inPKT[964]      = 112'hC2C47573206574206E6574757320;
        inPKT[965]      = 112'hC2C56574206D616C657375616461;
        inPKT[966]      = 112'hC2C62066616D6573206163207475;
        inPKT[967]      = 112'hC2C7727069732065676573746173;
        inPKT[968]      = 112'hC2C82E20496E206665726D656E74;
        inPKT[969]      = 112'hC2C9756D2061742075726E61206E;
        inPKT[970]      = 112'hC2CA6F6E20636F6E76616C6C6973;
        inPKT[971]      = 112'hC2CB2E20446F6E65632061632061;
        inPKT[972]      = 112'hC2CC75677565206A7573746F2E20;
        inPKT[973]      = 112'hC2CD496E20617420656C69742065;
        inPKT[974]      = 112'hC2CE742061726375206D6178696D;
        inPKT[975]      = 112'hC2CF7573206C75637475732E2046;
        inPKT[976]      = 112'hC2D07573636520657569736D6F64;
        inPKT[977]      = 112'hC2D1206E756E63206E6563207665;
        inPKT[978]      = 112'hC2D26E656E617469732061756374;
        inPKT[979]      = 112'hC2D36F722E204C6F72656D206970;
        inPKT[980]      = 112'hC2D473756D20646F6C6F72207369;
        inPKT[981]      = 112'hC2D57420616D65742C20636F6E73;
        inPKT[982]      = 112'hC2D6656374657475722061646970;
        inPKT[983]      = 112'hC2D7697363696E6720656C69742E;
        inPKT[984]      = 112'hC2D820446F6E6563206469637475;
        inPKT[985]      = 112'hC2D96D2074656D706F7220727574;
        inPKT[986]      = 112'hC2DA72756D2E2053656420656C65;
        inPKT[987]      = 112'hC2DB6966656E64206469616D2069;
        inPKT[988]      = 112'hC2DC64206D6173736120696D7065;
        inPKT[989]      = 112'hC2DD72646965742C206163206F72;
        inPKT[990]      = 112'hC2DE6E617265206C696265726F20;
        inPKT[991]      = 112'hC2DF656C656966656E642E204D61;
        inPKT[992]      = 112'hC2E06563656E6173206F726E6172;
        inPKT[993]      = 112'hC2E165206D65747573206E756C6C;
        inPKT[994]      = 112'hC2E2612C2073697420616D657420;
        inPKT[995]      = 112'hC2E36665726D656E74756D20656C;
        inPKT[996]      = 112'hC2E4697420616C697175616D2069;
        inPKT[997]      = 112'hC2E5642E20446F6E656320756C74;
        inPKT[998]      = 112'hC2E6726963657320746F72746F72;
        inPKT[999]      = 112'hC2E720617420616E74652068656E;
        inPKT[1000]     = 112'hC2E86472657269742C2065752073;
        inPKT[1001]     = 112'hC2E961676974746973206A757374;
        inPKT[1002]     = 112'hC2EA6F20756C7472696365732E0D;
        inPKT[1003]     = 112'hC2EB0A0D0A5072616573656E7420;
        inPKT[1004]     = 112'hC2EC6C7563747573207072657469;
        inPKT[1005]     = 112'hC2ED756D206E657175652C207369;
        inPKT[1006]     = 112'hC2EE7420616D65742070656C6C65;
        inPKT[1007]     = 112'hC2EF6E746573717565206D617572;
        inPKT[1008]     = 112'hC2F0697320656C656D656E74756D;
        inPKT[1009]     = 112'hC2F1206E6F6E2E20557420626C61;
        inPKT[1010]     = 112'hC2F26E6469742070686172657472;
        inPKT[1011]     = 112'hC2F361206F64696F206E6F6E2065;
        inPKT[1012]     = 112'hC2F47569736D6F642E2051756973;
        inPKT[1013]     = 112'hC2F5717565207669746165206C65;
        inPKT[1014]     = 112'hC2F66F20616C697175616D2C2073;
        inPKT[1015]     = 112'hC2F76F64616C65732074656C6C75;
        inPKT[1016]     = 112'hC2F8732069642C20696163756C69;
        inPKT[1017]     = 112'hC2F973206D61757269732E204E61;
        inPKT[1018]     = 112'hC2FA6D2065666669636974757220;
        inPKT[1019]     = 112'hC2FB696E20707572757320736564;
        inPKT[1020]     = 112'hC2FC20616363756D73616E2E204D;
        inPKT[1021]     = 112'hC2FD616563656E61732073697420;
        inPKT[1022]     = 112'hC2FE616D65742063757273757320;
        inPKT[1023]     = 112'hC2FF66656C69732E205175697371;
        inPKT[1024]     = 112'hC20075652066617563696275732C;
        inPKT[1025]     = 112'hC201206475692065742061756374;
        inPKT[1026]     = 112'hC2026F72206C75637475732C2061;
        inPKT[1027]     = 112'hC2036E7465206572617420706F73;
        inPKT[1028]     = 112'hC204756572652065726F732C2075;
        inPKT[1029]     = 112'hC2057420636F6E76616C6C697320;
        inPKT[1030]     = 112'hC2066D65747573206C6563747573;
        inPKT[1031]     = 112'hC207207669746165206C656F2E20;
        inPKT[1032]     = 112'hC20853757370656E646973736520;
        inPKT[1033]     = 112'hC209706F74656E74692E20437261;
        inPKT[1034]     = 112'hC20A7320657420646F6C6F72206E;
        inPKT[1035]     = 112'hC20B6F6E2075726E61207363656C;
        inPKT[1036]     = 112'hC20C657269737175652074726973;
        inPKT[1037]     = 112'hC20D74697175652E204372617320;
        inPKT[1038]     = 112'hC20E72757472756D206E65632076;
        inPKT[1039]     = 112'hC20F656C69742061632073616769;
        inPKT[1040]     = 112'hC210747469732E20446F6E656320;
        inPKT[1041]     = 112'hC211656C656966656E642C206C61;
        inPKT[1042]     = 112'hC212637573207365642067726176;
        inPKT[1043]     = 112'hC213696461206D616C6573756164;
        inPKT[1044]     = 112'hC214612C20657820616E74652070;
        inPKT[1045]     = 112'hC2156C616365726174206C656374;
        inPKT[1046]     = 112'hC21675732C206567657420636F6E;
        inPKT[1047]     = 112'hC217677565206D61737361206D65;
        inPKT[1048]     = 112'hC218747573206964206C61637573;
        inPKT[1049]     = 112'hC2192E2053757370656E64697373;
        inPKT[1050]     = 112'hC21A652069642072757472756D20;
        inPKT[1051]     = 112'hC21B6C65637475732E2046757363;
        inPKT[1052]     = 112'hC21C65206D6178696D7573207365;
        inPKT[1053]     = 112'hC21D64206C6967756C6120736564;
        inPKT[1054]     = 112'hC21E20766976657272612E204E61;
        inPKT[1055]     = 112'hC21F6D206C756374757320646961;
        inPKT[1056]     = 112'hC2206D20616E74652C2076697461;
        inPKT[1057]     = 112'hC22165206F726E617265206E6571;
        inPKT[1058]     = 112'hC222756520766172697573206567;
        inPKT[1059]     = 112'hC22365742E0D0A0D0A50656C6C65;
        inPKT[1060]     = 112'hC2246E7465737175652061742065;
        inPKT[1061]     = 112'hC2256C6974206E6962682E205665;
        inPKT[1062]     = 112'hC22673746962756C756D20616E74;
        inPKT[1063]     = 112'hC2276520697073756D207072696D;
        inPKT[1064]     = 112'hC228697320696E20666175636962;
        inPKT[1065]     = 112'hC2297573206F726369206C756374;
        inPKT[1066]     = 112'hC22A757320657420756C74726963;
        inPKT[1067]     = 112'hC22B657320706F73756572652063;
        inPKT[1068]     = 112'hC22C7562696C6961204375726165;
        inPKT[1069]     = 112'hC22D3B2043757261626974757220;
        inPKT[1070]     = 112'hC22E666175636962757320646961;
        inPKT[1071]     = 112'hC22F6D206C656F2C206E65632065;
        inPKT[1072]     = 112'hC2307569736D6F642073656D2065;
        inPKT[1073]     = 112'hC23166666963697475722075742E;
        inPKT[1074]     = 112'hC232205574207665686963756C61;
        inPKT[1075]     = 112'hC233206175677565206163206C69;
        inPKT[1076]     = 112'hC2346265726F20696163756C6973;
        inPKT[1077]     = 112'hC2352C206E656320656C65696665;
        inPKT[1078]     = 112'hC2366E6420657820706F7274612E;
        inPKT[1079]     = 112'hC237204D6F7262692068656E6472;
        inPKT[1080]     = 112'hC238657269742067726176696461;
        inPKT[1081]     = 112'hC2392074696E636964756E742E20;
        inPKT[1082]     = 112'hC23A5072616573656E7420646F6C;
        inPKT[1083]     = 112'hC23B6F72206C616375732C207465;
        inPKT[1084]     = 112'hC23C6D707573206575206672696E;
        inPKT[1085]     = 112'hC23D67696C6C612073697420616D;
        inPKT[1086]     = 112'hC23E65742C20656C656966656E64;
        inPKT[1087]     = 112'hC23F20696E206E756C6C612E204E;
        inPKT[1088]     = 112'hC240756C6C61206D6F6C6C697320;
        inPKT[1089]     = 112'hC24165676574206D61676E61206E;
        inPKT[1090]     = 112'hC24265632068656E647265726974;
        inPKT[1091]     = 112'hC2432E20416C697175616D20636F;
        inPKT[1092]     = 112'hC2446E76616C6C69732073656D20;
        inPKT[1093]     = 112'hC24576697461652073617069656E;
        inPKT[1094]     = 112'hC2462064696374756D2C20757420;
        inPKT[1095]     = 112'hC247766573746962756C756D206C;
        inPKT[1096]     = 112'hC2486F72656D206672696E67696C;
        inPKT[1097]     = 112'hC2496C612E20446F6E6563207465;
        inPKT[1098]     = 112'hC24A6C6C7573206C696265726F2C;
        inPKT[1099]     = 112'hC24B206665756769617420757420;
        inPKT[1100]     = 112'hC24C66696E69627573206E65632C;
        inPKT[1101]     = 112'hC24D20616C697175616D20736974;
        inPKT[1102]     = 112'hC24E20616D6574206F7263692E20;
        inPKT[1103]     = 112'hC24F4E756E632073757363697069;
        inPKT[1104]     = 112'hC25074206E69736C206574206F72;
        inPKT[1105]     = 112'hC2516E6172652076657374696275;
        inPKT[1106]     = 112'hC2526C756D2E204E756C6C616D20;
        inPKT[1107]     = 112'hC2536C6F626F7274697320736170;
        inPKT[1108]     = 112'hC25469656E206A7573746F2C2073;
        inPKT[1109]     = 112'hC255697420616D6574206469676E;
        inPKT[1110]     = 112'hC256697373696D206E756C6C6120;
        inPKT[1111]     = 112'hC257636F6E64696D656E74756D20;
        inPKT[1112]     = 112'hC258696E2E20536564206D6F6C65;
        inPKT[1113]     = 112'hC2597374696520766F6C75747061;
        inPKT[1114]     = 112'hC25A74206E697369206174206665;
        inPKT[1115]     = 112'hC25B726D656E74756D2E204E756C;
        inPKT[1116]     = 112'hC25C6C61206D6F6C657374696520;
        inPKT[1117]     = 112'hC25D6E6973692073656420747572;
        inPKT[1118]     = 112'hC25E706973206D6F6C6573746965;
        inPKT[1119]     = 112'hC25F2C206E6F6E20696163756C69;
        inPKT[1120]     = 112'hC26073206E756E63206661756369;
        inPKT[1121]     = 112'hC2616275732E2041656E65616E20;
        inPKT[1122]     = 112'hC262696E74657264756D20706861;
        inPKT[1123]     = 112'hC263726574726120636F6E736563;
        inPKT[1124]     = 112'hC26474657475722E20457469616D;
        inPKT[1125]     = 112'hC265206578206F7263692C206961;
        inPKT[1126]     = 112'hC26663756C6973206E6F6E206575;
        inPKT[1127]     = 112'hC26769736D6F642069642C20756C;
        inPKT[1128]     = 112'hC2686C616D636F72706572207363;
        inPKT[1129]     = 112'hC269656C65726973717565206F64;
        inPKT[1130]     = 112'hC26A696F2E0D0A0D0A4E616D2075;
        inPKT[1131]     = 112'hC26B6C74726963657320656C6569;
        inPKT[1132]     = 112'hC26C66656E64206469616D2C2065;
        inPKT[1133]     = 112'hC26D67657420736F64616C657320;
        inPKT[1134]     = 112'hC26E73656D206D61747469732061;
        inPKT[1135]     = 112'hC26F632E2055742076656E656E61;
        inPKT[1136]     = 112'hC270746973206E69626820657520;
        inPKT[1137]     = 112'hC2716C65637475732074696E6369;
        inPKT[1138]     = 112'hC27264756E742064696374756D2E;
        inPKT[1139]     = 112'hC27320566976616D757320637572;
        inPKT[1140]     = 112'hC274737573206175677565207175;
        inPKT[1141]     = 112'hC2756973206C6F626F7274697320;
        inPKT[1142]     = 112'hC276657569736D6F642E204E756E;
        inPKT[1143]     = 112'hC2776320616C697175616D206469;
        inPKT[1144]     = 112'hC278616D20617420616E74652066;
        inPKT[1145]     = 112'hC2796163696C69736973206D6178;
        inPKT[1146]     = 112'hC27A696D75732E20457469616D20;
        inPKT[1147]     = 112'hC27B736564206C6F72656D206D61;
        inPKT[1148]     = 112'hC27C747469732C20636F6E76616C;
        inPKT[1149]     = 112'hC27D6C69732075726E6120766974;
        inPKT[1150]     = 112'hC27E61652C2074656D7075732073;
        inPKT[1151]     = 112'hC27F656D2E20566976616D757320;
        inPKT[1152]     = 112'hC2806567657374617320766F6C75;
        inPKT[1153]     = 112'hC281747061742065726F73206575;
        inPKT[1154]     = 112'hC28220756C7472696365732E2056;
        inPKT[1155]     = 112'hC2836573746962756C756D20756C;
        inPKT[1156]     = 112'hC2846C616D636F72706572206572;
        inPKT[1157]     = 112'hC2856174206E756E632C206E6F6E;
        inPKT[1158]     = 112'hC2862068656E647265726974206F;
        inPKT[1159]     = 112'hC28764696F2070656C6C656E7465;
        inPKT[1160]     = 112'hC288737175652069642E20467573;
        inPKT[1161]     = 112'hC28963652075726E612069707375;
        inPKT[1162]     = 112'hC28A6D2C206C6163696E69612069;
        inPKT[1163]     = 112'hC28B6E2073757363697069742076;
        inPKT[1164]     = 112'hC28C656C2C2073656D7065722069;
        inPKT[1165]     = 112'hC28D6E206F64696F2E2050656C6C;
        inPKT[1166]     = 112'hC28E656E74657371756520696420;
        inPKT[1167]     = 112'hC28F6E696268206E6973692E2041;
        inPKT[1168]     = 112'hC2906C697175616D20706F727461;
        inPKT[1169]     = 112'hC291206E69736C20657420657820;
        inPKT[1170]     = 112'hC292696163756C69732074726973;
        inPKT[1171]     = 112'hC29374697175652E20457469616D;
        inPKT[1172]     = 112'hC294206D61737361206F7263692C;
        inPKT[1173]     = 112'hC295206567657374617320736564;
        inPKT[1174]     = 112'hC296206C6F72656D20717569732C;
        inPKT[1175]     = 112'hC297206469676E697373696D2073;
        inPKT[1176]     = 112'hC298656D70657220616E74652E20;
        inPKT[1177]     = 112'hC29953757370656E646973736520;
        inPKT[1178]     = 112'hC29A74696E636964756E74206E69;
        inPKT[1179]     = 112'hC29B73692065782C207365642076;
        inPKT[1180]     = 112'hC29C6F6C75747061742065737420;
        inPKT[1181]     = 112'hC29D766172697573207669746165;
        inPKT[1182]     = 112'hC29E2E0D0A0D0A5365642073656D;
        inPKT[1183]     = 112'hC29F706572206C6163696E696120;
        inPKT[1184]     = 112'hC2A0646F6C6F722E204E616D2075;
        inPKT[1185]     = 112'hC2A1742076656C697420696E206C;
        inPKT[1186]     = 112'hC2A26163757320636F6E73656374;
        inPKT[1187]     = 112'hC2A36574757220636F6E76616C6C;
        inPKT[1188]     = 112'hC2A469732070656C6C656E746573;
        inPKT[1189]     = 112'hC2A5717565207365642073656D2E;
        inPKT[1190]     = 112'hC2A62053757370656E6469737365;
        inPKT[1191]     = 112'hC2A720636F6E64696D656E74756D;
        inPKT[1192]     = 112'hC2A820612065726F732069642075;
        inPKT[1193]     = 112'hC2A96C6C616D636F727065722E20;
        inPKT[1194]     = 112'hC2AA4D6F726269206C7563747573;
        inPKT[1195]     = 112'hC2AB2075726E612073697420616D;
        inPKT[1196]     = 112'hC2AC657420657569736D6F642069;
        inPKT[1197]     = 112'hC2AD6163756C69732E2050656C6C;
        inPKT[1198]     = 112'hC2AE656E74657371756520666163;
        inPKT[1199]     = 112'hC2AF696C69736973206D61757269;
        inPKT[1200]     = 112'hC2B07320657520656C656D656E74;
        inPKT[1201]     = 112'hC2B1756D207661726975732E204F;
        inPKT[1202]     = 112'hC2B272636920766172697573206E;
        inPKT[1203]     = 112'hC2B361746F7175652070656E6174;
        inPKT[1204]     = 112'hC2B469627573206574206D61676E;
        inPKT[1205]     = 112'hC2B5697320646973207061727475;
        inPKT[1206]     = 112'hC2B67269656E74206D6F6E746573;
        inPKT[1207]     = 112'hC2B72C206E617363657475722072;
        inPKT[1208]     = 112'hC2B869646963756C7573206D7573;
        inPKT[1209]     = 112'hC2B92E20446F6E6563206469676E;
        inPKT[1210]     = 112'hC2BA697373696D20612069707375;
        inPKT[1211]     = 112'hC2BB6D20756C7472696369657320;
        inPKT[1212]     = 112'hC2BC76656E656E617469732E2056;
        inPKT[1213]     = 112'hC2BD6976616D7573206E756E6320;
        inPKT[1214]     = 112'hC2BE76656C69742C207665686963;
        inPKT[1215]     = 112'hC2BF756C61207669746165206D61;
        inPKT[1216]     = 112'hC2C07373612075742C20636F6E76;
        inPKT[1217]     = 112'hC2C1616C6C697320636F6E736563;
        inPKT[1218]     = 112'hC2C2746574757220746F72746F72;
        inPKT[1219]     = 112'hC2C32E205175697371756520616C;
        inPKT[1220]     = 112'hC2C4697175616D2C206E69736C20;
        inPKT[1221]     = 112'hC2C5636F6E67756520626C616E64;
        inPKT[1222]     = 112'hC2C6697420756C74726963696573;
        inPKT[1223]     = 112'hC2C72C2075726E61207475727069;
        inPKT[1224]     = 112'hC2C873206D6174746973206D6167;
        inPKT[1225]     = 112'hC2C96E612C206E6F6E206665726D;
        inPKT[1226]     = 112'hC2CA656E74756D20647569207665;
        inPKT[1227]     = 112'hC2CB6C6974206575207175616D2E;
        inPKT[1228]     = 112'hC2CC0D0A0D0A496E207068617265;
        inPKT[1229]     = 112'hC2CD7472612076656C697420646F;
        inPKT[1230]     = 112'hC2CE6C6F722C2076697461652063;
        inPKT[1231]     = 112'hC2CF7572737573206F7263692066;
        inPKT[1232]     = 112'hC2D0696E696275732074696E6369;
        inPKT[1233]     = 112'hC2D164756E742E20566976616D75;
        inPKT[1234]     = 112'hC2D27320696420746F72746F7220;
        inPKT[1235]     = 112'hC2D372686F6E6375732C20736167;
        inPKT[1236]     = 112'hC2D46974746973206469616D2065;
        inPKT[1237]     = 112'hC2D56765742C207072657469756D;
        inPKT[1238]     = 112'hC2D6206D61757269732E20506861;
        inPKT[1239]     = 112'hC2D773656C6C757320656C656D65;
        inPKT[1240]     = 112'hC2D86E74756D20656E696D206665;
        inPKT[1241]     = 112'hC2D96C69732E204D617572697320;
        inPKT[1242]     = 112'hC2DA6575206E6571756520656765;
        inPKT[1243]     = 112'hC2DB742070757275732068656E64;
        inPKT[1244]     = 112'hC2DC726572697420677261766964;
        inPKT[1245]     = 112'hC2DD612E20416C697175616D206C;
        inPKT[1246]     = 112'hC2DE696265726F206E6962682C20;
        inPKT[1247]     = 112'hC2DF636F6E76616C6C6973206120;
        inPKT[1248]     = 112'hC2E06E69736C2065742C2068656E;
        inPKT[1249]     = 112'hC2E1647265726974207665737469;
        inPKT[1250]     = 112'hC2E262756C756D2066656C69732E;
        inPKT[1251]     = 112'hC2E320446F6E656320657569736D;
        inPKT[1252]     = 112'hC2E46F64206665726D656E74756D;
        inPKT[1253]     = 112'hC2E5207475727069732065752061;
        inPKT[1254]     = 112'hC2E67563746F722E2041656E6561;
        inPKT[1255]     = 112'hC2E76E20626962656E64756D2074;
        inPKT[1256]     = 112'hC2E8757270697320696E206F6469;
        inPKT[1257]     = 112'hC2E96F20636F6E76616C6C69732C;
        inPKT[1258]     = 112'hC2EA207669746165207661726975;
        inPKT[1259]     = 112'hC2EB73206578206C616F72656574;
        inPKT[1260]     = 112'hC2EC2E2046757363652076656C20;
        inPKT[1261]     = 112'hC2ED6D6920766974616520646F6C;
        inPKT[1262]     = 112'hC2EE6F7220666575676961742076;
        inPKT[1263]     = 112'hC2EF756C707574617465206E6563;
        inPKT[1264]     = 112'hC2F0207574206E756E632E204372;
        inPKT[1265]     = 112'hC2F1617320646170696275732C20;
        inPKT[1266]     = 112'hC2F2616E74652069642076656869;
        inPKT[1267]     = 112'hC2F363756C6120616C697175616D;
        inPKT[1268]     = 112'hC2F42C20656C69742065726F7320;
        inPKT[1269]     = 112'hC2F57361676974746973206D692C;
        inPKT[1270]     = 112'hC2F6206E6F6E20656C656966656E;
        inPKT[1271]     = 112'hC2F764206578206E756C6C612065;
        inPKT[1272]     = 112'hC2F86765742076656C69742E2053;
        inPKT[1273]     = 112'hC2F9757370656E64697373652069;
        inPKT[1274]     = 112'hC2FA64206469616D206475692E20;
        inPKT[1275]     = 112'hC2FB53757370656E646973736520;
        inPKT[1276]     = 112'hC2FC7072657469756D206A757374;
        inPKT[1277]     = 112'hC2FD6F20736564206E6962682070;
        inPKT[1278]     = 112'hC2FE6F72747469746F722C207665;
        inPKT[1279]     = 112'hC2FF6C20696E74657264756D206D;
        inPKT[1280]     = 112'hC2006175726973206D6178696D75;
        inPKT[1281]     = 112'hC201732E20557420616C69717561;
        inPKT[1282]     = 112'hC2026D206C616375732070757275;
        inPKT[1283]     = 112'hC203732C2073697420616D657420;
        inPKT[1284]     = 112'hC204696D70657264696574206E69;
        inPKT[1285]     = 112'hC205626820666575676961742069;
        inPKT[1286]     = 112'hC206642E20496E7465676572206C;
        inPKT[1287]     = 112'hC2076F72656D206D61757269732C;
        inPKT[1288]     = 112'hC208207072657469756D206E6F6E;
        inPKT[1289]     = 112'hC209206E6973692065742C206461;
        inPKT[1290]     = 112'hC20A70696275732066696E696275;
        inPKT[1291]     = 112'hC20B73206F7263692E0D0A0D0A56;
        inPKT[1292]     = 112'hC20C6573746962756C756D206961;
        inPKT[1293]     = 112'hC20D63756C69732C206D61676E61;
        inPKT[1294]     = 112'hC20E206174206D6174746973206D;
        inPKT[1295]     = 112'hC20F6178696D75732C2061726375;
        inPKT[1296]     = 112'hC210206572617420646170696275;
        inPKT[1297]     = 112'hC21173206E756E632C2061207661;
        inPKT[1298]     = 112'hC21272697573206D657475732066;
        inPKT[1299]     = 112'hC213656C697320736564206F7263;
        inPKT[1300]     = 112'hC214692E204E756C6C616D206D69;
        inPKT[1301]     = 112'hC215206E6962682C20656C656966;
        inPKT[1302]     = 112'hC216656E64206E656320756C7472;
        inPKT[1303]     = 112'hC21769636573206E65632C20636F;
        inPKT[1304]     = 112'hC2186E7365637465747572206163;
        inPKT[1305]     = 112'hC21920656E696D2E20536564206C;
        inPKT[1306]     = 112'hC21A75637475732073656D207175;
        inPKT[1307]     = 112'hC21B69732074656D706F7220636F;
        inPKT[1308]     = 112'hC21C6E6775652E2053757370656E;
        inPKT[1309]     = 112'hC21D646973736520706F74656E74;
        inPKT[1310]     = 112'hC21E692E20457469616D20656765;
        inPKT[1311]     = 112'hC21F74206C696265726F2076656C;
        inPKT[1312]     = 112'hC22069742E204475697320766573;
        inPKT[1313]     = 112'hC221746962756C756D20636F6E73;
        inPKT[1314]     = 112'hC222657175617420706F7274612E;
        inPKT[1315]     = 112'hC223204D617572697320706F7274;
        inPKT[1316]     = 112'hC2247469746F7220747572706973;
        inPKT[1317]     = 112'hC22520696E206D6173736120616C;
        inPKT[1318]     = 112'hC226697175616D20636F6E677565;
        inPKT[1319]     = 112'hC2272E204E756C6C6120636F6E73;
        inPKT[1320]     = 112'hC228656374657475722075726E61;
        inPKT[1321]     = 112'hC229206D657475732C2069642069;
        inPKT[1322]     = 112'hC22A6163756C6973206E756E6320;
        inPKT[1323]     = 112'hC22B756C74726963696573206567;
        inPKT[1324]     = 112'hC22C65742E204375726162697475;
        inPKT[1325]     = 112'hC22D72206D6175726973206E6571;
        inPKT[1326]     = 112'hC22E75652C20626962656E64756D;
        inPKT[1327]     = 112'hC22F207365642065726F73206174;
        inPKT[1328]     = 112'hC2302C206D6178696D757320756C;
        inPKT[1329]     = 112'hC231747269636573207475727069;
        inPKT[1330]     = 112'hC232732E0D0A496E74657264756D;
        inPKT[1331]     = 112'hC233206574206D616C6573756164;
        inPKT[1332]     = 112'hC234612066616D65732061632061;
        inPKT[1333]     = 112'hC2356E746520697073756D207072;
        inPKT[1334]     = 112'hC236696D697320696E2066617563;
        inPKT[1335]     = 112'hC237696275732E2050656C6C656E;
        inPKT[1336]     = 112'hC23874657371756520736F6C6C69;
        inPKT[1337]     = 112'hC2396369747564696E20626C616E;
        inPKT[1338]     = 112'hC23A646974206665726D656E7475;
        inPKT[1339]     = 112'hC23B6D2E2050656C6C656E746573;
        inPKT[1340]     = 112'hC23C717565206E6F6E206C696775;
        inPKT[1341]     = 112'hC23D6C6120657520657261742076;
        inPKT[1342]     = 112'hC23E656E656E6174697320657569;
        inPKT[1343]     = 112'hC23F736D6F642E2050656C6C656E;
        inPKT[1344]     = 112'hC24074657371756520736F64616C;
        inPKT[1345]     = 112'hC241657320766573746962756C75;
        inPKT[1346]     = 112'hC2426D20636F6E76616C6C69732E;
        inPKT[1347]     = 112'hC2432050726F696E206D6F6C6573;
        inPKT[1348]     = 112'hC244746965207072657469756D20;
        inPKT[1349]     = 112'hC24565726F732076656C20656765;
        inPKT[1350]     = 112'hC246737461732E204D6F72626920;
        inPKT[1351]     = 112'hC247736F6C6C696369747564696E;
        inPKT[1352]     = 112'hC248207075727573206163206665;
        inPKT[1353]     = 112'hC249726D656E74756D206D617474;
        inPKT[1354]     = 112'hC24A69732E204E756E632076656C;
        inPKT[1355]     = 112'hC24B2074696E636964756E74206C;
        inPKT[1356]     = 112'hC24C696265726F2E204E756C6C61;
        inPKT[1357]     = 112'hC24D20616C697175657420697073;
        inPKT[1358]     = 112'hC24E756D206E6563207175616D20;
        inPKT[1359]     = 112'hC24F696D7065726469657420696E;
        inPKT[1360]     = 112'hC25074657264756D2E2050726165;
        inPKT[1361]     = 112'hC25173656E74206C6967756C6120;
        inPKT[1362]     = 112'hC25266656C69732C20696163756C;
        inPKT[1363]     = 112'hC253697320617420616C69717565;
        inPKT[1364]     = 112'hC254742061742C20736167697474;
        inPKT[1365]     = 112'hC2556973207175697320656C6974;
        inPKT[1366]     = 112'hC2562E0D0A517569737175652076;
        inPKT[1367]     = 112'hC257656C20696D70657264696574;
        inPKT[1368]     = 112'hC258206E6962682E205068617365;
        inPKT[1369]     = 112'hC2596C6C75732072757472756D20;
        inPKT[1370]     = 112'hC25A6469676E697373696D207269;
        inPKT[1371]     = 112'hC25B737573206E6F6E2074696E63;
        inPKT[1372]     = 112'hC25C6964756E742E205665737469;
        inPKT[1373]     = 112'hC25D62756C756D206E756E632069;
        inPKT[1374]     = 112'hC25E7073756D2C2076656E656E61;
        inPKT[1375]     = 112'hC25F746973206567657420706F72;
        inPKT[1376]     = 112'hC260746120696E2C20636F6E7365;
        inPKT[1377]     = 112'hC261637465747572206575206572;
        inPKT[1378]     = 112'hC26261742E20446F6E6563207665;
        inPKT[1379]     = 112'hC263686963756C6120616E746520;
        inPKT[1380]     = 112'hC26476656C2072686F6E63757320;
        inPKT[1381]     = 112'hC26566617563696275732E205065;
        inPKT[1382]     = 112'hC2666C6C656E746573717565206A;
        inPKT[1383]     = 112'hC2677573746F20746F72746F722C;
        inPKT[1384]     = 112'hC26820766F6C757470617420696E;
        inPKT[1385]     = 112'hC269206D61757269732061742C20;
        inPKT[1386]     = 112'hC26A766172697573207068617265;
        inPKT[1387]     = 112'hC26B7472612072697375732E2051;
        inPKT[1388]     = 112'hC26C756973717565207574206469;
        inPKT[1389]     = 112'hC26D616D2073757363697069742C;
        inPKT[1390]     = 112'hC26E20736F6C6C69636974756469;
        inPKT[1391]     = 112'hC26F6E2073617069656E2065742C;
        inPKT[1392]     = 112'hC27020696E74657264756D206C61;
        inPKT[1393]     = 112'hC2716375732E204D6F7262692072;
        inPKT[1394]     = 112'hC272697375732073656D2C207065;
        inPKT[1395]     = 112'hC2736C6C656E7465737175652065;
        inPKT[1396]     = 112'hC274742074757270697320696E2C;
        inPKT[1397]     = 112'hC27520626C616E64697420736F6C;
        inPKT[1398]     = 112'hC2766C696369747564696E207365;
        inPKT[1399]     = 112'hC2776D2E20536564206566666963;
        inPKT[1400]     = 112'hC27869747572206C696265726F20;
        inPKT[1401]     = 112'hC27971756973207072657469756D;
        inPKT[1402]     = 112'hC27A207072657469756D2E204E75;
        inPKT[1403]     = 112'hC27B6C6C616D20617563746F7220;
        inPKT[1404]     = 112'hC27C7361676974746973206C6F72;
        inPKT[1405]     = 112'hC27D656D2C20616320756C747269;
        inPKT[1406]     = 112'hC27E6365732061726375206D6178;
        inPKT[1407]     = 112'hC27F696D757320656765742E0D0A;
        inPKT[1408]     = 112'hC280566573746962756C756D2076;
        inPKT[1409]     = 112'hC2816F6C7574706174206C696775;
        inPKT[1410]     = 112'hC2826C6120617563746F72207365;
        inPKT[1411]     = 112'hC2836D20766976657272612C2075;
        inPKT[1412]     = 112'hC2846C6C616D636F727065722065;
        inPKT[1413]     = 112'hC2857569736D6F64206E65717565;
        inPKT[1414]     = 112'hC28620706F72747469746F722E20;
        inPKT[1415]     = 112'hC28753757370656E646973736520;
        inPKT[1416]     = 112'hC28876697665727261207363656C;
        inPKT[1417]     = 112'hC28965726973717565206F64696F;
        inPKT[1418]     = 112'hC28A2072686F6E63757320766F6C;
        inPKT[1419]     = 112'hC28B75747061742E20416C697175;
        inPKT[1420]     = 112'hC28C616D206572617420766F6C75;
        inPKT[1421]     = 112'hC28D747061742E2053757370656E;
        inPKT[1422]     = 112'hC28E646973736520706F74656E74;
        inPKT[1423]     = 112'hC28F692E20496E20686163206861;
        inPKT[1424]     = 112'hC2906269746173736520706C6174;
        inPKT[1425]     = 112'hC29165612064696374756D73742E;
        inPKT[1426]     = 112'hC2922050726F696E207574206E75;
        inPKT[1427]     = 112'hC2936C6C61207574206475692073;
        inPKT[1428]     = 112'hC29463656C657269737175652064;
        inPKT[1429]     = 112'hC295696374756D2E205175697371;
        inPKT[1430]     = 112'hC296756520737573636970697420;
        inPKT[1431]     = 112'hC2976E69626820706F7375657265;
        inPKT[1432]     = 112'hC298207175616D2076756C707574;
        inPKT[1433]     = 112'hC2996174652C206575206C616369;
        inPKT[1434]     = 112'hC29A6E696120616E746520677261;
        inPKT[1435]     = 112'hC29B766964612E20437572616269;
        inPKT[1436]     = 112'hC29C747572206D61737361206C6F;
        inPKT[1437]     = 112'hC29D72656D2C206F726E61726520;
        inPKT[1438]     = 112'hC29E6575206D6F6C6C6973206174;
        inPKT[1439]     = 112'hC29F2C207068617265747261206E;
        inPKT[1440]     = 112'hC2A06563206D617373612E204E75;
        inPKT[1441]     = 112'hC2A16C6C612066696E6962757320;
        inPKT[1442]     = 112'hC2A2656C656966656E64206F7263;
        inPKT[1443]     = 112'hC2A3692073697420616D65742063;
        inPKT[1444]     = 112'hC2A46F6E73656374657475722E20;
        inPKT[1445]     = 112'hC2A55365642074656D7075732076;
        inPKT[1446]     = 112'hC2A6697461652061726375206E65;
        inPKT[1447]     = 112'hC2A763206665726D656E74756D2E;
        inPKT[1448]     = 112'hC2A82041656E65616E2070656C6C;
        inPKT[1449]     = 112'hC2A9656E74657371756520766974;
        inPKT[1450]     = 112'hC2AA616520646F6C6F7220696E20;
        inPKT[1451]     = 112'hC2AB616363756D73616E2E204372;
        inPKT[1452]     = 112'hC2AC6173206469676E697373696D;
        inPKT[1453]     = 112'hC2AD2076756C707574617465206D;
        inPKT[1454]     = 112'hC2AE6F6C6C69732E204D61757269;
        inPKT[1455]     = 112'hC2AF7320706F7274612076656E65;
        inPKT[1456]     = 112'hC2B06E617469732072697375732C;
        inPKT[1457]     = 112'hC2B1206575207472697374697175;
        inPKT[1458]     = 112'hC2B26520646F6C6F722072757472;
        inPKT[1459]     = 112'hC2B3756D20696E2E204675736365;
        inPKT[1460]     = 112'hC2B420636F6E64696D656E74756D;
        inPKT[1461]     = 112'hC2B5206F7263692066656C69732C;
        inPKT[1462]     = 112'hC2B62073697420616D657420636F;
        inPKT[1463]     = 112'hC2B76E76616C6C6973206C696265;
        inPKT[1464]     = 112'hC2B8726F2074696E636964756E74;
        inPKT[1465]     = 112'hC2B92061632E0D0A566573746962;
        inPKT[1466]     = 112'hC2BA756C756D20696D7065726469;
        inPKT[1467]     = 112'hC2BB657420656C69742074656D70;
        inPKT[1468]     = 112'hC2BC6F72207175616D2067726176;
        inPKT[1469]     = 112'hC2BD6964612C207574206D616C65;
        inPKT[1470]     = 112'hC2BE73756164612074656C6C7573;
        inPKT[1471]     = 112'hC2BF20696D706572646965742E20;
        inPKT[1472]     = 112'hC2C050686173656C6C7573206F64;
        inPKT[1473]     = 112'hC2C1696F2073656D2C206D617474;
        inPKT[1474]     = 112'hC2C269732073656420756C747269;
        inPKT[1475]     = 112'hC2C36365732061742C2076697665;
        inPKT[1476]     = 112'hC2C47272612076656C206475692E;
        inPKT[1477]     = 112'hC2C5204E756E632075726E61206D;
        inPKT[1478]     = 112'hC2C6657475732C206C7563747573;
        inPKT[1479]     = 112'hC2C7206163206D6178696D757320;
        inPKT[1480]     = 112'hC2C8696E2C20636F6E7365637465;
        inPKT[1481]     = 112'hC2C9747572206E6F6E206E697369;
        inPKT[1482]     = 112'hC2CA2E204E756C6C612073697420;
        inPKT[1483]     = 112'hC2CB616D657420626962656E6475;
        inPKT[1484]     = 112'hC2CC6D2076656C69742E20446F6E;
        inPKT[1485]     = 112'hC2CD6563207175697320656E696D;
        inPKT[1486]     = 112'hC2CE206E6F6E2072697375732062;
        inPKT[1487]     = 112'hC2CF6C616E64697420666163696C;
        inPKT[1488]     = 112'hC2D0697369732071756973206E65;
        inPKT[1489]     = 112'hC2D1632072697375732E20437572;
        inPKT[1490]     = 112'hC2D2616269747572206575206573;
        inPKT[1491]     = 112'hC2D374207669746165206C656374;
        inPKT[1492]     = 112'hC2D4757320626C616E6469742061;
        inPKT[1493]     = 112'hC2D56C69717565742E2056657374;
        inPKT[1494]     = 112'hC2D66962756C756D20616E746520;
        inPKT[1495]     = 112'hC2D7697073756D207072696D6973;
        inPKT[1496]     = 112'hC2D820696E206661756369627573;
        inPKT[1497]     = 112'hC2D9206F726369206C7563747573;
        inPKT[1498]     = 112'hC2DA20657420756C747269636573;
        inPKT[1499]     = 112'hC2DB20706F737565726520637562;
        inPKT[1500]     = 112'hC2DC696C69612043757261653B20;
        inPKT[1501]     = 112'hC2DD566573746962756C756D2061;
        inPKT[1502]     = 112'hC2DE63206469676E697373696D20;
        inPKT[1503]     = 112'hC2DF6E756E632E20517569737175;
        inPKT[1504]     = 112'hC2E06520696E2073616769747469;
        inPKT[1505]     = 112'hC2E1732074656C6C75732C207369;
        inPKT[1506]     = 112'hC2E27420616D6574206665726D65;
        inPKT[1507]     = 112'hC2E36E74756D206E6962682E0D0A;
        inPKT[1508]     = 112'hC2E4496E206469676E697373696D;
        inPKT[1509]     = 112'hC2E5207269737573207669746165;
        inPKT[1510]     = 112'hC2E6207075727573207665737469;
        inPKT[1511]     = 112'hC2E762756C756D2C20617420656C;
        inPKT[1512]     = 112'hC2E8656D656E74756D206E756C6C;
        inPKT[1513]     = 112'hC2E96120706F73756572652E2053;
        inPKT[1514]     = 112'hC2EA6564206D6174746973206E75;
        inPKT[1515]     = 112'hC2EB6E63206E6962682E20537573;
        inPKT[1516]     = 112'hC2EC70656E64697373652070656C;
        inPKT[1517]     = 112'hC2ED6C656E74657371756520706C;
        inPKT[1518]     = 112'hC2EE616365726174207363656C65;
        inPKT[1519]     = 112'hC2EF7269737175652E2041656E65;
        inPKT[1520]     = 112'hC2F0616E2066657567696174206D;
        inPKT[1521]     = 112'hC2F1617572697320696420636F6E;
        inPKT[1522]     = 112'hC2F2677565206C6163696E69612E;
        inPKT[1523]     = 112'hC2F320457469616D207375736369;
        inPKT[1524]     = 112'hC2F4706974206C6967756C612074;
        inPKT[1525]     = 112'hC2F5656C6C75732C206120636F6E;
        inPKT[1526]     = 112'hC2F6677565206C65637475732061;
        inPKT[1527]     = 112'hC2F76C697175616D207665686963;
        inPKT[1528]     = 112'hC2F8756C612E2053757370656E64;
        inPKT[1529]     = 112'hC2F969737365206567657420616E;
        inPKT[1530]     = 112'hC2FA74652076656C20656E696D20;
        inPKT[1531]     = 112'hC2FB6D616C657375616461207669;
        inPKT[1532]     = 112'hC2FC76657272612E2050726F696E;
        inPKT[1533]     = 112'hC2FD2074696E636964756E742061;
        inPKT[1534]     = 112'hC2FE72637520656765742076756C;
        inPKT[1535]     = 112'hC2FF70757461746520616363756D;
        inPKT[1536]     = 112'hC20073616E2E20496E2076697461;
        inPKT[1537]     = 112'hC20165206469616D206E6962682E;
        inPKT[1538]     = 112'hC202204D6F726269206D6178696D;
        inPKT[1539]     = 112'hC20375732066656C697320696420;
        inPKT[1540]     = 112'hC204636F6E736563746574757220;
        inPKT[1541]     = 112'hC205616C697175616D2E204E756C;
        inPKT[1542]     = 112'hC2066C6120666163696C6973692E;
        inPKT[1543]     = 112'hC2070D0A566573746962756C756D;
        inPKT[1544]     = 112'hC20820766573746962756C756D20;
        inPKT[1545]     = 112'hC20965666669636974757220746F;
        inPKT[1546]     = 112'hC20A72746F722073697420616D65;
        inPKT[1547]     = 112'hC20B7420666163696C697369732E;
        inPKT[1548]     = 112'hC20C204D616563656E6173206E6F;
        inPKT[1549]     = 112'hC20D6E2074656C6C7573206F7263;
        inPKT[1550]     = 112'hC20E692E2050686173656C6C7573;
        inPKT[1551]     = 112'hC20F206E6F6E206C756374757320;
        inPKT[1552]     = 112'hC2106A7573746F2C206174207375;
        inPKT[1553]     = 112'hC2117363697069742074656C6C75;
        inPKT[1554]     = 112'hC212732E2046757363652068656E;
        inPKT[1555]     = 112'hC213647265726974206E6563206E;
        inPKT[1556]     = 112'hC2146962682076656C2063757273;
        inPKT[1557]     = 112'hC21575732E2053757370656E6469;
        inPKT[1558]     = 112'hC21673736520706F74656E74692E;
        inPKT[1559]     = 112'hC2172044756973206C6967756C61;
        inPKT[1560]     = 112'hC2182066656C69732C2065666669;
        inPKT[1561]     = 112'hC21963697475722065742076656C;
        inPKT[1562]     = 112'hC21A69742061742C20666163696C;
        inPKT[1563]     = 112'hC21B6973697320636F6E76616C6C;
        inPKT[1564]     = 112'hC21C6973206A7573746F2E204E75;
        inPKT[1565]     = 112'hC21D6C6C616D206C6F626F727469;
        inPKT[1566]     = 112'hC21E732070656C6C656E74657371;
        inPKT[1567]     = 112'hC21F756520736F6C6C6963697475;
        inPKT[1568]     = 112'hC22064696E2E204E616D20736974;
        inPKT[1569]     = 112'hC22120616D657420646F6C6F7220;
        inPKT[1570]     = 112'hC22273697420616D6574206C6563;
        inPKT[1571]     = 112'hC22374757320696D706572646965;
        inPKT[1572]     = 112'hC2247420636F6E7365717561742E;
        inPKT[1573]     = 112'hC22520416C697175616D206C7563;
        inPKT[1574]     = 112'hC226747573207363656C65726973;
        inPKT[1575]     = 112'hC2277175652070757275732C2069;
        inPKT[1576]     = 112'hC22864206672696E67696C6C6120;
        inPKT[1577]     = 112'hC22973656D20766F6C7574706174;
        inPKT[1578]     = 112'hC22A2061632E205365642074656D;
        inPKT[1579]     = 112'hC22B706F722C20656E696D206567;
        inPKT[1580]     = 112'hC22C657420657569736D6F642066;
        inPKT[1581]     = 112'hC22D6163696C697369732C206E69;
        inPKT[1582]     = 112'hC22E73692065782073656D706572;
        inPKT[1583]     = 112'hC22F20697073756D2C20696E2073;
        inPKT[1584]     = 112'hC23061676974746973206F726369;
        inPKT[1585]     = 112'hC231207175616D20696E206C6563;
        inPKT[1586]     = 112'hC2327475732E2055742076697461;
        inPKT[1587]     = 112'hC2336520656C6974206C6967756C;
        inPKT[1588]     = 112'hC234612E204E756E632065676573;
        inPKT[1589]     = 112'hC2357461732C206D692076697461;
        inPKT[1590]     = 112'hC2366520696163756C6973206D61;
        inPKT[1591]     = 112'hC237747469732C20647569206E69;
        inPKT[1592]     = 112'hC238626820656C656966656E6420;
        inPKT[1593]     = 112'hC2396E69736C2C20656765742070;
        inPKT[1594]     = 112'hC23A6F727461206C696265726F20;
        inPKT[1595]     = 112'hC23B617567756520717569732065;
        inPKT[1596]     = 112'hC23C6E696D2E2053656420736974;
        inPKT[1597]     = 112'hC23D20616D65742070756C76696E;
        inPKT[1598]     = 112'hC23E61722065782C2076656C2070;
        inPKT[1599]     = 112'hC23F656C6C656E74657371756520;
        inPKT[1600]     = 112'hC2406C61637573206E756C6C616D;

	in = inPKT[countIN];

	@(posedge clk);
	#10ns

	nR = 1'b1;

	@(posedge clk);
	#10ns
	
	in_newPKT <= 1'b1;
end

always @(posedge clk)				countCYCLE <= countCYCLE + 1'b1;

always @(posedge in_loadPKT)
begin
	repeat(2)	@(posedge clk);
	#10ns
	
	if(~doneSIM && (countIN != `PKT_MAX))	countIN <= countIN + 1'b1;
	else					doneSIM = 1'b1;
	in_newPKT <= 1'b0;
end

always @(posedge in_donePKT)
begin
	repeat(2)	@(posedge clk);
	#10ns

	if(~doneSIM)
	begin
		in = inPKT[countIN];
	
		@(posedge clk)
		in_newPKT <= 1'b1;
	end
end

always @(posedge out_donePKT)
begin
	if(countOUT != `PKT_MAX)		countOUT <= countOUT + 1'b1;
	else
	begin
		$display("%d PACKETS PROCESS AND FINISHED @ %tns in %d cycles", countOUT, $time, countCYCLE);
	end

	repeat(2)	@(posedge clk);
	#10ns
	
	out_readPKT <= 1'b1;

	repeat(2)	@(posedge clk);
	#10ns

	out_readPKT <= 1'b0;
end

endmodule
